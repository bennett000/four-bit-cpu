.title KiCad schematic
.tran 1ns 2000ns
.print tran v(Din) v(ClkIn) v(ClrIn) v(CEIn) v(flipflopdclrceQ)
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V1 flipflopdclrceVcc 0 dc 5
V2 Din 0 dc 5
V3 ClkIn 0 PULSE(0 5 2NS 2NS 2NS 50NS 100NS)
V4 ClrIn 0 dc 5
V5 CEIn 0 dc 0
R3 flipflopdclrceVcc flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor2A 1K
R1 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
R2 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
Q1 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor2A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1AorB 0 NPN
R6 flipflopdclrceVcc flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3A 1K
R4 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor2A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
R5 flipflopdclrceCEandClk flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
Q2 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor2AorB 0 NPN
R10 flipflopdclrceVcc flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4A 1K
R7 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R8 flipflopdclrceCEandClk flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
Q3 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 0 NPN
R9 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R13 flipflopdclrceVcc flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1A 1K
R11 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
R12 Din flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
Q4 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor1A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4AorB 0 NPN
R17 flipflopdclrceVcc flipflopdclrceQ 1K
R14 ClrIn flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R15 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor3A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
Q5 flipflopdclrceQ flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 0 NPN
R16 flipflopdclrceNQ flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R20 flipflopdclrceVcc flipflopdclrceNQ 1K
R18 flipflopdclrceQ flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
R19 flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor4A flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
Q6 flipflopdclrceNQ flipflopdclrceflipflopdclrceflipflopdclrflipflopdclrnor6AorB 0 NPN
R23 flipflopdclrceVcc flipflopdclrceCEandClk 1K
R21 flipflopdclrceflipflopdclrceand1sheet5C364DB7A flipflopdclrceflipflopdclrceand1sheet5C364DB7AorB 10K
R22 flipflopdclrceflipflopdclrceand1sheet5C364DB7B flipflopdclrceflipflopdclrceand1sheet5C364DB7AorB 10K
Q7 flipflopdclrceCEandClk flipflopdclrceflipflopdclrceand1sheet5C364DB7AorB 0 NPN
R25 flipflopdclrceVcc flipflopdclrceflipflopdclrceand1sheet5C364DB7A 1K
R24 ClkIn flipflopdclrceflipflopdclrceand1Sheet5C3654CCQr 10K
Q8 flipflopdclrceflipflopdclrceand1sheet5C364DB7A flipflopdclrceflipflopdclrceand1Sheet5C3654CCQr 0 NPN
R27 flipflopdclrceVcc flipflopdclrceflipflopdclrceand1sheet5C364DB7B 1K
R26 CEIn flipflopdclrceflipflopdclrceand1sheet5C366192Qr 10K
Q9 flipflopdclrceflipflopdclrceand1sheet5C364DB7B flipflopdclrceflipflopdclrceand1sheet5C366192Qr 0 NPN
.end
