.title KiCad schematic
.tran 1ns 2000ns
.print tran v(ClkIn) v(ClrIn) v(CEIn) v(register4q1) v(register4q2) v(register4q3) v(register4q4)
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V2 register4Vcc 0 dc 5
V1 D1In 0 dc 5
V6 ClkIn 0 PULSE(0 5 2NS 2NS 2NS 50NS 100NS)
V7 ClrIn 0 dc 0
V8 CEIn 0 dc 5
V3 D2In 0 dc 0
V4 D3In 0 dc 5
V5 D4In 0 dc 5
R3 register4Vcc register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor2A 1K
R1 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
R2 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
Q1 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1AorB 0 NPN
R6 register4Vcc register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3A 1K
R4 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
R5 register4register4flipflop1CEandClk register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
Q2 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor2AorB 0 NPN
R10 register4Vcc register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4A 1K
R7 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R8 register4register4flipflop1CEandClk register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
Q3 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 0 NPN
R9 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R13 register4Vcc register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1A 1K
R11 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
R12 D1In register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
Q4 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4AorB 0 NPN
R17 register4Vcc register4Q1 1K
R14 ClrIn register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R15 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
Q5 register4Q1 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 0 NPN
R16 register4NQ1 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R20 register4Vcc register4NQ1 1K
R18 register4Q1 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
R19 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
Q6 register4NQ1 register4register4flipflop1flipflopdclrceflipflopdclrflipflopdclrnor6AorB 0 NPN
R23 register4Vcc register4register4flipflop1CEandClk 1K
R21 register4register4flipflop1flipflopdclrceand1sheet5C364DB7A register4register4flipflop1flipflopdclrceand1sheet5C364DB7AorB 10K
R22 register4register4flipflop1flipflopdclrceand1sheet5C364DB7B register4register4flipflop1flipflopdclrceand1sheet5C364DB7AorB 10K
Q7 register4register4flipflop1CEandClk register4register4flipflop1flipflopdclrceand1sheet5C364DB7AorB 0 NPN
R25 register4Vcc register4register4flipflop1flipflopdclrceand1sheet5C364DB7A 1K
R24 ClkIn register4register4flipflop1flipflopdclrceand1Sheet5C3654CCQr 10K
Q8 register4register4flipflop1flipflopdclrceand1sheet5C364DB7A register4register4flipflop1flipflopdclrceand1Sheet5C3654CCQr 0 NPN
R27 register4Vcc register4register4flipflop1flipflopdclrceand1sheet5C364DB7B 1K
R26 CEIn register4register4flipflop1flipflopdclrceand1sheet5C366192Qr 10K
Q9 register4register4flipflop1flipflopdclrceand1sheet5C364DB7B register4register4flipflop1flipflopdclrceand1sheet5C366192Qr 0 NPN
R30 register4Vcc register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor2A 1K
R28 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
R29 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
Q10 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1AorB 0 NPN
R33 register4Vcc register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3A 1K
R31 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
R32 register4register4flipflop2CEandClk register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
Q11 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor2AorB 0 NPN
R37 register4Vcc register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4A 1K
R34 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R35 register4register4flipflop2CEandClk register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
Q12 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 0 NPN
R36 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R40 register4Vcc register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1A 1K
R38 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
R39 D2In register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
Q13 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4AorB 0 NPN
R44 register4Vcc register4Q2 1K
R41 ClrIn register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R42 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
Q14 register4Q2 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 0 NPN
R43 register4NQ2 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R47 register4Vcc register4NQ2 1K
R45 register4Q2 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
R46 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
Q15 register4NQ2 register4register4flipflop2flipflopdclrceflipflopdclrflipflopdclrnor6AorB 0 NPN
R50 register4Vcc register4register4flipflop2CEandClk 1K
R48 register4register4flipflop2flipflopdclrceand1sheet5C364DB7A register4register4flipflop2flipflopdclrceand1sheet5C364DB7AorB 10K
R49 register4register4flipflop2flipflopdclrceand1sheet5C364DB7B register4register4flipflop2flipflopdclrceand1sheet5C364DB7AorB 10K
Q16 register4register4flipflop2CEandClk register4register4flipflop2flipflopdclrceand1sheet5C364DB7AorB 0 NPN
R52 register4Vcc register4register4flipflop2flipflopdclrceand1sheet5C364DB7A 1K
R51 ClkIn register4register4flipflop2flipflopdclrceand1Sheet5C3654CCQr 10K
Q17 register4register4flipflop2flipflopdclrceand1sheet5C364DB7A register4register4flipflop2flipflopdclrceand1Sheet5C3654CCQr 0 NPN
R54 register4Vcc register4register4flipflop2flipflopdclrceand1sheet5C364DB7B 1K
R53 CEIn register4register4flipflop2flipflopdclrceand1sheet5C366192Qr 10K
Q18 register4register4flipflop2flipflopdclrceand1sheet5C364DB7B register4register4flipflop2flipflopdclrceand1sheet5C366192Qr 0 NPN
R57 register4Vcc register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor2A 1K
R55 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
R56 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
Q19 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1AorB 0 NPN
R60 register4Vcc register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3A 1K
R58 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
R59 register4register4flipflop3CEandClk register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
Q20 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor2AorB 0 NPN
R64 register4Vcc register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4A 1K
R61 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R62 register4register4flipflop3CEandClk register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
Q21 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 0 NPN
R63 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R67 register4Vcc register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1A 1K
R65 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
R66 D3In register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
Q22 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4AorB 0 NPN
R71 register4Vcc register4Q3 1K
R68 ClrIn register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R69 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
Q23 register4Q3 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 0 NPN
R70 register4NQ3 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R74 register4Vcc register4NQ3 1K
R72 register4Q3 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
R73 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
Q24 register4NQ3 register4register4flipflop3flipflopdclrceflipflopdclrflipflopdclrnor6AorB 0 NPN
R77 register4Vcc register4register4flipflop3CEandClk 1K
R75 register4register4flipflop3flipflopdclrceand1sheet5C364DB7A register4register4flipflop3flipflopdclrceand1sheet5C364DB7AorB 10K
R76 register4register4flipflop3flipflopdclrceand1sheet5C364DB7B register4register4flipflop3flipflopdclrceand1sheet5C364DB7AorB 10K
Q25 register4register4flipflop3CEandClk register4register4flipflop3flipflopdclrceand1sheet5C364DB7AorB 0 NPN
R79 register4Vcc register4register4flipflop3flipflopdclrceand1sheet5C364DB7A 1K
R78 ClkIn register4register4flipflop3flipflopdclrceand1Sheet5C3654CCQr 10K
Q26 register4register4flipflop3flipflopdclrceand1sheet5C364DB7A register4register4flipflop3flipflopdclrceand1Sheet5C3654CCQr 0 NPN
R81 register4Vcc register4register4flipflop3flipflopdclrceand1sheet5C364DB7B 1K
R80 CEIn register4register4flipflop3flipflopdclrceand1sheet5C366192Qr 10K
Q27 register4register4flipflop3flipflopdclrceand1sheet5C364DB7B register4register4flipflop3flipflopdclrceand1sheet5C366192Qr 0 NPN
R84 register4Vcc register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor2A 1K
R82 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
R83 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1AorB 10K
Q28 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1AorB 0 NPN
R87 register4Vcc register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3A 1K
R85 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor2A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
R86 register4register4flipflop4CEandClk register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor2AorB 10K
Q29 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor2AorB 0 NPN
R91 register4Vcc register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4A 1K
R88 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R89 register4register4flipflop4CEandClk register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
Q30 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 0 NPN
R90 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3AorBorC 10K
R94 register4Vcc register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1A 1K
R92 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
R93 D4In register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4AorB 10K
Q31 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor1A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4AorB 0 NPN
R98 register4Vcc register4Q4 1K
R95 ClrIn register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R96 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor3A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
Q32 register4Q4 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 0 NPN
R97 register4NQ4 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor5AorBorC 10K
R101 register4Vcc register4NQ4 1K
R99 register4Q4 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
R100 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor4A register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor6AorB 10K
Q33 register4NQ4 register4register4flipflop4flipflopdclrceflipflopdclrflipflopdclrnor6AorB 0 NPN
R104 register4Vcc register4register4flipflop4CEandClk 1K
R102 register4register4flipflop4flipflopdclrceand1sheet5C364DB7A register4register4flipflop4flipflopdclrceand1sheet5C364DB7AorB 10K
R103 register4register4flipflop4flipflopdclrceand1sheet5C364DB7B register4register4flipflop4flipflopdclrceand1sheet5C364DB7AorB 10K
Q34 register4register4flipflop4CEandClk register4register4flipflop4flipflopdclrceand1sheet5C364DB7AorB 0 NPN
R106 register4Vcc register4register4flipflop4flipflopdclrceand1sheet5C364DB7A 1K
R105 ClkIn register4register4flipflop4flipflopdclrceand1Sheet5C3654CCQr 10K
Q35 register4register4flipflop4flipflopdclrceand1sheet5C364DB7A register4register4flipflop4flipflopdclrceand1Sheet5C3654CCQr 0 NPN
R108 register4Vcc register4register4flipflop4flipflopdclrceand1sheet5C364DB7B 1K
R107 CEIn register4register4flipflop4flipflopdclrceand1sheet5C366192Qr 10K
Q36 register4register4flipflop4flipflopdclrceand1sheet5C364DB7B register4register4flipflop4flipflopdclrceand1sheet5C366192Qr 0 NPN
.end
