.title KiCad schematic
.op
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V2 bitwiseinv44Vcc 0 dc 5
V1 En 0 dc 5
V3 A1 0 dc 5
V4 A2 0 dc 0
V5 A3 0 dc 5
V6 A4 0 dc 0
R3 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor21xor2nor2B 1K
R1 En bitwiseinv44bitwiseinvxor21xor2nor1AorB 10K
R2 A1 bitwiseinv44bitwiseinvxor21xor2nor1AorB 10K
Q1 bitwiseinv44bitwiseinvxor21xor2nor2B bitwiseinv44bitwiseinvxor21xor2nor1AorB 0 NPN
R6 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor21xor2nor2A 1K
R4 bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7AorB 10K
R5 bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7AorB 10K
Q2 bitwiseinv44bitwiseinvxor21xor2nor2A bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7AorB 0 NPN
R8 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7A 1K
R7 En bitwiseinv44bitwiseinvxor21xor2and1Sheet5C3654CCQr 10K
Q3 bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor21xor2and1Sheet5C3654CCQr 0 NPN
R10 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7B 1K
R9 A1 bitwiseinv44bitwiseinvxor21xor2and1sheet5C366192Qr 10K
Q4 bitwiseinv44bitwiseinvxor21xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor21xor2and1sheet5C366192Qr 0 NPN
R13 bitwiseinv44Vcc bitwiseinv44Z1 1K
R11 bitwiseinv44bitwiseinvxor21xor2nor2A bitwiseinv44bitwiseinvxor21xor2nor2AorB 10K
R12 bitwiseinv44bitwiseinvxor21xor2nor2B bitwiseinv44bitwiseinvxor21xor2nor2AorB 10K
Q5 bitwiseinv44Z1 bitwiseinv44bitwiseinvxor21xor2nor2AorB 0 NPN
R16 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor22xor2nor2B 1K
R14 En bitwiseinv44bitwiseinvxor22xor2nor1AorB 10K
R15 A2 bitwiseinv44bitwiseinvxor22xor2nor1AorB 10K
Q6 bitwiseinv44bitwiseinvxor22xor2nor2B bitwiseinv44bitwiseinvxor22xor2nor1AorB 0 NPN
R19 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor22xor2nor2A 1K
R17 bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7AorB 10K
R18 bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7AorB 10K
Q7 bitwiseinv44bitwiseinvxor22xor2nor2A bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7AorB 0 NPN
R21 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7A 1K
R20 En bitwiseinv44bitwiseinvxor22xor2and1Sheet5C3654CCQr 10K
Q8 bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor22xor2and1Sheet5C3654CCQr 0 NPN
R23 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7B 1K
R22 A2 bitwiseinv44bitwiseinvxor22xor2and1sheet5C366192Qr 10K
Q9 bitwiseinv44bitwiseinvxor22xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor22xor2and1sheet5C366192Qr 0 NPN
R26 bitwiseinv44Vcc bitwiseinv44Z2 1K
R24 bitwiseinv44bitwiseinvxor22xor2nor2A bitwiseinv44bitwiseinvxor22xor2nor2AorB 10K
R25 bitwiseinv44bitwiseinvxor22xor2nor2B bitwiseinv44bitwiseinvxor22xor2nor2AorB 10K
Q10 bitwiseinv44Z2 bitwiseinv44bitwiseinvxor22xor2nor2AorB 0 NPN
R29 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor23xor2nor2B 1K
R27 En bitwiseinv44bitwiseinvxor23xor2nor1AorB 10K
R28 A3 bitwiseinv44bitwiseinvxor23xor2nor1AorB 10K
Q11 bitwiseinv44bitwiseinvxor23xor2nor2B bitwiseinv44bitwiseinvxor23xor2nor1AorB 0 NPN
R32 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor23xor2nor2A 1K
R30 bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7AorB 10K
R31 bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7AorB 10K
Q12 bitwiseinv44bitwiseinvxor23xor2nor2A bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7AorB 0 NPN
R34 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7A 1K
R33 En bitwiseinv44bitwiseinvxor23xor2and1Sheet5C3654CCQr 10K
Q13 bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor23xor2and1Sheet5C3654CCQr 0 NPN
R36 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7B 1K
R35 A3 bitwiseinv44bitwiseinvxor23xor2and1sheet5C366192Qr 10K
Q14 bitwiseinv44bitwiseinvxor23xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor23xor2and1sheet5C366192Qr 0 NPN
R39 bitwiseinv44Vcc bitwiseinv44Z3 1K
R37 bitwiseinv44bitwiseinvxor23xor2nor2A bitwiseinv44bitwiseinvxor23xor2nor2AorB 10K
R38 bitwiseinv44bitwiseinvxor23xor2nor2B bitwiseinv44bitwiseinvxor23xor2nor2AorB 10K
Q15 bitwiseinv44Z3 bitwiseinv44bitwiseinvxor23xor2nor2AorB 0 NPN
R42 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor24xor2nor2B 1K
R40 En bitwiseinv44bitwiseinvxor24xor2nor1AorB 10K
R41 A4 bitwiseinv44bitwiseinvxor24xor2nor1AorB 10K
Q16 bitwiseinv44bitwiseinvxor24xor2nor2B bitwiseinv44bitwiseinvxor24xor2nor1AorB 0 NPN
R45 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor24xor2nor2A 1K
R43 bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7AorB 10K
R44 bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7AorB 10K
Q17 bitwiseinv44bitwiseinvxor24xor2nor2A bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7AorB 0 NPN
R47 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7A 1K
R46 En bitwiseinv44bitwiseinvxor24xor2and1Sheet5C3654CCQr 10K
Q18 bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7A bitwiseinv44bitwiseinvxor24xor2and1Sheet5C3654CCQr 0 NPN
R49 bitwiseinv44Vcc bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7B 1K
R48 A4 bitwiseinv44bitwiseinvxor24xor2and1sheet5C366192Qr 10K
Q19 bitwiseinv44bitwiseinvxor24xor2and1sheet5C364DB7B bitwiseinv44bitwiseinvxor24xor2and1sheet5C366192Qr 0 NPN
R52 bitwiseinv44Vcc bitwiseinv44Z4 1K
R50 bitwiseinv44bitwiseinvxor24xor2nor2A bitwiseinv44bitwiseinvxor24xor2nor2AorB 10K
R51 bitwiseinv44bitwiseinvxor24xor2nor2B bitwiseinv44bitwiseinvxor24xor2nor2AorB 10K
Q20 bitwiseinv44Z4 bitwiseinv44bitwiseinvxor24xor2nor2AorB 0 NPN
.end
