.title KiCad schematic
V1 /and-2/Vcc 0 dc 5
V2 /Ain 0 dc 5
V3 /Bin 0 dc 5
R3 /and-2/Vcc /Q 1K
R1 /and-2/sheet5C364DB7/A /and-2/sheet5C364DB7/AorB 10K
R2 /and-2/sheet5C364DB7/B /and-2/sheet5C364DB7/AorB 10K
Q1 /Q /and-2/sheet5C364DB7/AorB 0 NPN
R5 /and-2/Vcc /and-2/sheet5C364DB7/A 1K
R4 /Ain /and-2/Sheet5C3654CC/Qr 10K
Q2 /and-2/sheet5C364DB7/A /and-2/Sheet5C3654CC/Qr 0 NPN
R7 /and-2/Vcc /and-2/sheet5C364DB7/B 1K
R6 /Bin /and-2/sheet5C366192/Qr 10K
Q3 /and-2/sheet5C364DB7/B /and-2/sheet5C366192/Qr 0 NPN
.end
