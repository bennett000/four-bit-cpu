.title KiCad schematic
.op
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V1 multiplexer441Vcc 0 dc 5
V2 A1in 0 dc 5
V3 A2in 0 dc 0
V4 A3in 0 dc 0
V5 A4in 0 dc 0
V9 B4in 0 dc 0
V8 B3in 0 dc 0
V7 B2in 0 dc 5
V6 B1in 0 dc 0
V18 multiplexer441S1 0 dc 5
V13 C4in 0 dc 0
V12 C3in 0 dc 0
V11 C2in 0 dc 5
V10 C1in 0 dc 5
V17 D4in 0 dc 0
V16 D3in 0 dc 5
V15 D2in 0 dc 0
V14 D1in 0 dc 0
V19 multiplexer441S2 0 dc 5
R2 multiplexer441Vcc multiplexer441multiplexer441mux4213A1 1K
R1 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornot1Qr 10K
Q1 multiplexer441multiplexer441mux4213A1 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R5 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornor1Q 1K
R3 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornor1AorB 10K
R4 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornor1AorB 10K
Q2 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R8 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1A 1K
R6 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R7 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q3 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R10 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R9 A1in multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q4 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R12 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R11 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q5 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R15 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1B 1K
R13 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R14 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q6 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R17 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R16 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q7 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R19 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R18 B1in multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q8 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R21 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1B 1K
R20 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21not1Qr 10K
Q9 multiplexer441multiplexer441mux4211multiplexer421mux1211mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1211mux21not1Qr 0 NPN
R23 multiplexer441Vcc multiplexer441multiplexer441mux4213A2 1K
R22 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornot1Qr 10K
Q10 multiplexer441multiplexer441mux4213A2 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R26 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornor1Q 1K
R24 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornor1AorB 10K
R25 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornor1AorB 10K
Q11 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R29 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1A 1K
R27 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R28 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q12 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R31 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R30 A2in multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q13 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R33 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R32 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q14 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R36 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1B 1K
R34 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R35 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q15 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R38 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R37 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q16 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R40 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R39 B2in multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q17 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R42 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1B 1K
R41 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21not1Qr 10K
Q18 multiplexer441multiplexer441mux4211multiplexer421mux1212mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1212mux21not1Qr 0 NPN
R44 multiplexer441Vcc multiplexer441multiplexer441mux4213A3 1K
R43 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornot1Qr 10K
Q19 multiplexer441multiplexer441mux4213A3 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R47 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornor1Q 1K
R45 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornor1AorB 10K
R46 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornor1AorB 10K
Q20 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R50 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1A 1K
R48 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R49 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q21 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R52 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R51 A3in multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q22 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R54 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R53 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q23 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R57 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1B 1K
R55 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R56 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q24 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R59 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R58 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q25 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R61 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R60 B3in multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q26 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R63 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1B 1K
R62 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21not1Qr 10K
Q27 multiplexer441multiplexer441mux4211multiplexer421mux1213mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1213mux21not1Qr 0 NPN
R65 multiplexer441Vcc multiplexer441multiplexer441mux4213A4 1K
R64 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornot1Qr 10K
Q28 multiplexer441multiplexer441mux4213A4 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R68 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornor1Q 1K
R66 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornor1AorB 10K
R67 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornor1AorB 10K
Q29 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornor1Q multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R71 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1A 1K
R69 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R70 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q30 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1A multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R73 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R72 A4in multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q31 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R75 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R74 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q32 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R78 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1B 1K
R76 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R77 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q33 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21or1B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R80 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R79 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q34 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R82 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R81 B4in multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q35 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R84 multiplexer441Vcc multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1B 1K
R83 multiplexer441S1 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21not1Qr 10K
Q36 multiplexer441multiplexer441mux4211multiplexer421mux1214mux21and1B multiplexer441multiplexer441mux4211multiplexer421mux1214mux21not1Qr 0 NPN
R86 multiplexer441Vcc multiplexer441multiplexer441mux4213B1 1K
R85 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornot1Qr 10K
Q37 multiplexer441multiplexer441mux4213B1 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R89 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornor1Q 1K
R87 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornor1AorB 10K
R88 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornor1AorB 10K
Q38 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R92 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1A 1K
R90 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R91 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q39 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R94 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R93 C1in multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q40 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R96 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R95 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q41 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R99 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1B 1K
R97 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R98 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q42 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R101 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R100 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q43 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R103 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R102 D1in multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q44 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R105 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1B 1K
R104 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21not1Qr 10K
Q45 multiplexer441multiplexer441mux4212multiplexer421mux1211mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1211mux21not1Qr 0 NPN
R107 multiplexer441Vcc multiplexer441multiplexer441mux4213B2 1K
R106 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornot1Qr 10K
Q46 multiplexer441multiplexer441mux4213B2 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R110 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornor1Q 1K
R108 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornor1AorB 10K
R109 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornor1AorB 10K
Q47 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R113 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1A 1K
R111 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R112 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q48 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R115 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R114 C2in multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q49 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R117 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R116 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q50 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R120 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1B 1K
R118 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R119 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q51 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R122 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R121 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q52 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R124 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R123 D2in multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q53 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R126 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1B 1K
R125 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21not1Qr 10K
Q54 multiplexer441multiplexer441mux4212multiplexer421mux1212mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1212mux21not1Qr 0 NPN
R128 multiplexer441Vcc multiplexer441multiplexer441mux4213B3 1K
R127 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornot1Qr 10K
Q55 multiplexer441multiplexer441mux4213B3 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R131 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornor1Q 1K
R129 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornor1AorB 10K
R130 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornor1AorB 10K
Q56 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R134 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1A 1K
R132 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R133 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q57 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R136 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R135 C3in multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q58 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R138 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R137 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q59 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R141 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1B 1K
R139 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R140 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q60 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R143 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R142 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q61 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R145 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R144 D3in multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q62 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R147 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1B 1K
R146 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21not1Qr 10K
Q63 multiplexer441multiplexer441mux4212multiplexer421mux1213mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1213mux21not1Qr 0 NPN
R149 multiplexer441Vcc multiplexer441multiplexer441mux4213B4 1K
R148 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornot1Qr 10K
Q64 multiplexer441multiplexer441mux4213B4 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R152 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornor1Q 1K
R150 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornor1AorB 10K
R151 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornor1AorB 10K
Q65 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornor1Q multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R155 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1A 1K
R153 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R154 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q66 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1A multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R157 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R156 C4in multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q67 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R159 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R158 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q68 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R162 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1B 1K
R160 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R161 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q69 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21or1B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R164 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R163 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q70 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R166 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R165 D4in multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q71 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R168 multiplexer441Vcc multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1B 1K
R167 multiplexer441S1 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21not1Qr 10K
Q72 multiplexer441multiplexer441mux4212multiplexer421mux1214mux21and1B multiplexer441multiplexer441mux4212multiplexer421mux1214mux21not1Qr 0 NPN
R170 multiplexer441Vcc multiplexer441Z1 1K
R169 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornot1Qr 10K
Q73 multiplexer441Z1 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R173 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornor1Q 1K
R171 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornor1AorB 10K
R172 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornor1AorB 10K
Q74 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R176 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1A 1K
R174 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R175 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q75 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R178 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R177 multiplexer441multiplexer441mux4213A1 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q76 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R180 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R179 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q77 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R183 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1B 1K
R181 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R182 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q78 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R185 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R184 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q79 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R187 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R186 multiplexer441multiplexer441mux4213B1 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q80 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R189 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1B 1K
R188 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21not1Qr 10K
Q81 multiplexer441multiplexer441mux4213multiplexer421mux1211mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1211mux21not1Qr 0 NPN
R191 multiplexer441Vcc multiplexer441Z2 1K
R190 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornot1Qr 10K
Q82 multiplexer441Z2 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R194 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornor1Q 1K
R192 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornor1AorB 10K
R193 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornor1AorB 10K
Q83 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R197 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1A 1K
R195 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R196 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q84 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R199 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R198 multiplexer441multiplexer441mux4213A2 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q85 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R201 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R200 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q86 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R204 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1B 1K
R202 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R203 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q87 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R206 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R205 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q88 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R208 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R207 multiplexer441multiplexer441mux4213B2 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q89 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R210 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1B 1K
R209 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21not1Qr 10K
Q90 multiplexer441multiplexer441mux4213multiplexer421mux1212mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1212mux21not1Qr 0 NPN
R212 multiplexer441Vcc multiplexer441Z3 1K
R211 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornot1Qr 10K
Q91 multiplexer441Z3 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R215 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornor1Q 1K
R213 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornor1AorB 10K
R214 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornor1AorB 10K
Q92 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R218 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1A 1K
R216 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R217 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q93 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R220 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R219 multiplexer441multiplexer441mux4213A3 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q94 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R222 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R221 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q95 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R225 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1B 1K
R223 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R224 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q96 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R227 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R226 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q97 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R229 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R228 multiplexer441multiplexer441mux4213B3 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q98 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R231 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1B 1K
R230 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21not1Qr 10K
Q99 multiplexer441multiplexer441mux4213multiplexer421mux1213mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1213mux21not1Qr 0 NPN
R233 multiplexer441Vcc multiplexer441Z4 1K
R232 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornot1Qr 10K
Q100 multiplexer441Z4 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R236 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornor1Q 1K
R234 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornor1AorB 10K
R235 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornor1AorB 10K
Q101 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornor1Q multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R239 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1A 1K
R237 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R238 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q102 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1A multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R241 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R240 multiplexer441multiplexer441mux4213A4 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q103 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R243 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R242 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q104 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R246 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1B 1K
R244 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R245 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q105 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21or1B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R248 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R247 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q106 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R250 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R249 multiplexer441multiplexer441mux4213B4 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q107 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R252 multiplexer441Vcc multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1B 1K
R251 multiplexer441S2 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21not1Qr 10K
Q108 multiplexer441multiplexer441mux4213multiplexer421mux1214mux21and1B multiplexer441multiplexer441mux4213multiplexer421mux1214mux21not1Qr 0 NPN
.end
