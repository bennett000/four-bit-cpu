.model LED D (IS=1a RS=3.3 N=1.8)

