.title KiCad schematic
.model NPN npn (is=6.7e15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V1 adder4Vcc 0 dc -5
V4 register4aCLK 0 dc 0
V2 register4aD1 0 dc 0
V3 register4bD1 0 dc 0
R3 adder4Vcc adder4adder41sheet5C34B00DA 1K
R1 adder4A1 adder4adder41sheet5C34AF27AorB 10K
R2 adder4B1 adder4adder41sheet5C34AF27AorB 10K
Q1 adder4adder41sheet5C34B00DA adder4adder41sheet5C34AF27AorB 0 NPN
R6 adder4Vcc adder4adder41sheet5C34B027A 1K
R4 adder4A1 adder4adder41sheet5C34AFF9AorB 10K
R5 adder4adder41sheet5C34B00DA adder4adder41sheet5C34AFF9AorB 10K
Q2 adder4adder41sheet5C34B027A adder4adder41sheet5C34AFF9AorB 0 NPN
R9 adder4Vcc adder4adder41sheet5C34B027B 1K
R7 adder4adder41sheet5C34B00DA adder4adder41sheet5C34B00DAorB 10K
R8 adder4B1 adder4adder41sheet5C34B00DAorB 10K
Q3 adder4adder41sheet5C34B027B adder4adder41sheet5C34B00DAorB 0 NPN
R12 adder4Vcc adder4adder41sheet5C34B047A 1K
R10 adder4adder41sheet5C34B027A adder4adder41sheet5C34B027AorB 10K
R11 adder4adder41sheet5C34B027B adder4adder41sheet5C34B027AorB 10K
Q4 adder4adder41sheet5C34B047A adder4adder41sheet5C34B027AorB 0 NPN
R15 adder4Vcc adder4adder41sheet5C34B049A 1K
R13 adder4adder41sheet5C34B047A adder4adder41sheet5C34B047AorB 10K
R14 adder4Cin adder4adder41sheet5C34B047AorB 10K
Q5 adder4adder41sheet5C34B049A adder4adder41sheet5C34B047AorB 0 NPN
R18 adder4Vcc adder4adder41sheet5C34B04AA 1K
R16 adder4adder41sheet5C34B047A adder4adder41sheet5C34B048AorB 10K
R17 adder4adder41sheet5C34B049A adder4adder41sheet5C34B048AorB 10K
Q6 adder4adder41sheet5C34B04AA adder4adder41sheet5C34B048AorB 0 NPN
R21 adder4Vcc adder4adder41sheet5C34B04AB 1K
R19 adder4adder41sheet5C34B049A adder4adder41sheet5C34B049AorB 10K
R20 adder4Cin adder4adder41sheet5C34B049AorB 10K
Q7 adder4adder41sheet5C34B04AB adder4adder41sheet5C34B049AorB 0 NPN
R24 adder4Vcc register4rD1 1K
R22 adder4adder41sheet5C34B04AA adder4adder41sheet5C34B04AAorB 10K
R23 adder4adder41sheet5C34B04AB adder4adder41sheet5C34B04AAorB 10K
Q8 register4rD1 adder4adder41sheet5C34B04AAorB 0 NPN
R27 adder4Vcc adder4adder42Cin 1K
R25 adder4adder41sheet5C34B049A adder4adder41sheet5C34B0CDAorB 10K
R26 adder4adder41sheet5C34B00DA adder4adder41sheet5C34B0CDAorB 10K
Q9 adder4adder42Cin adder4adder41sheet5C34B0CDAorB 0 NPN
R30 adder4Vcc adder4adder42sheet5C34B00DA 1K
R28 adder4A2 adder4adder42sheet5C34AF27AorB 10K
R29 adder4B2 adder4adder42sheet5C34AF27AorB 10K
Q10 adder4adder42sheet5C34B00DA adder4adder42sheet5C34AF27AorB 0 NPN
R33 adder4Vcc adder4adder42sheet5C34B027A 1K
R31 adder4A2 adder4adder42sheet5C34AFF9AorB 10K
R32 adder4adder42sheet5C34B00DA adder4adder42sheet5C34AFF9AorB 10K
Q11 adder4adder42sheet5C34B027A adder4adder42sheet5C34AFF9AorB 0 NPN
R36 adder4Vcc adder4adder42sheet5C34B027B 1K
R34 adder4adder42sheet5C34B00DA adder4adder42sheet5C34B00DAorB 10K
R35 adder4B2 adder4adder42sheet5C34B00DAorB 10K
Q12 adder4adder42sheet5C34B027B adder4adder42sheet5C34B00DAorB 0 NPN
R39 adder4Vcc adder4adder42sheet5C34B047A 1K
R37 adder4adder42sheet5C34B027A adder4adder42sheet5C34B027AorB 10K
R38 adder4adder42sheet5C34B027B adder4adder42sheet5C34B027AorB 10K
Q13 adder4adder42sheet5C34B047A adder4adder42sheet5C34B027AorB 0 NPN
R42 adder4Vcc adder4adder42sheet5C34B049A 1K
R40 adder4adder42sheet5C34B047A adder4adder42sheet5C34B047AorB 10K
R41 adder4adder42Cin adder4adder42sheet5C34B047AorB 10K
Q14 adder4adder42sheet5C34B049A adder4adder42sheet5C34B047AorB 0 NPN
R45 adder4Vcc adder4adder42sheet5C34B04AA 1K
R43 adder4adder42sheet5C34B047A adder4adder42sheet5C34B048AorB 10K
R44 adder4adder42sheet5C34B049A adder4adder42sheet5C34B048AorB 10K
Q15 adder4adder42sheet5C34B04AA adder4adder42sheet5C34B048AorB 0 NPN
R48 adder4Vcc adder4adder42sheet5C34B04AB 1K
R46 adder4adder42sheet5C34B049A adder4adder42sheet5C34B049AorB 10K
R47 adder4adder42Cin adder4adder42sheet5C34B049AorB 10K
Q16 adder4adder42sheet5C34B04AB adder4adder42sheet5C34B049AorB 0 NPN
R51 adder4Vcc register4rD2 1K
R49 adder4adder42sheet5C34B04AA adder4adder42sheet5C34B04AAorB 10K
R50 adder4adder42sheet5C34B04AB adder4adder42sheet5C34B04AAorB 10K
Q17 register4rD2 adder4adder42sheet5C34B04AAorB 0 NPN
R54 adder4Vcc adder4adder43Cin 1K
R52 adder4adder42sheet5C34B049A adder4adder42sheet5C34B0CDAorB 10K
R53 adder4adder42sheet5C34B00DA adder4adder42sheet5C34B0CDAorB 10K
Q18 adder4adder43Cin adder4adder42sheet5C34B0CDAorB 0 NPN
R57 adder4Vcc adder4adder43sheet5C34B00DA 1K
R55 adder4A3 adder4adder43sheet5C34AF27AorB 10K
R56 adder4B3 adder4adder43sheet5C34AF27AorB 10K
Q19 adder4adder43sheet5C34B00DA adder4adder43sheet5C34AF27AorB 0 NPN
R60 adder4Vcc adder4adder43sheet5C34B027A 1K
R58 adder4A3 adder4adder43sheet5C34AFF9AorB 10K
R59 adder4adder43sheet5C34B00DA adder4adder43sheet5C34AFF9AorB 10K
Q20 adder4adder43sheet5C34B027A adder4adder43sheet5C34AFF9AorB 0 NPN
R63 adder4Vcc adder4adder43sheet5C34B027B 1K
R61 adder4adder43sheet5C34B00DA adder4adder43sheet5C34B00DAorB 10K
R62 adder4B3 adder4adder43sheet5C34B00DAorB 10K
Q21 adder4adder43sheet5C34B027B adder4adder43sheet5C34B00DAorB 0 NPN
R66 adder4Vcc adder4adder43sheet5C34B047A 1K
R64 adder4adder43sheet5C34B027A adder4adder43sheet5C34B027AorB 10K
R65 adder4adder43sheet5C34B027B adder4adder43sheet5C34B027AorB 10K
Q22 adder4adder43sheet5C34B047A adder4adder43sheet5C34B027AorB 0 NPN
R69 adder4Vcc adder4adder43sheet5C34B049A 1K
R67 adder4adder43sheet5C34B047A adder4adder43sheet5C34B047AorB 10K
R68 adder4adder43Cin adder4adder43sheet5C34B047AorB 10K
Q23 adder4adder43sheet5C34B049A adder4adder43sheet5C34B047AorB 0 NPN
R72 adder4Vcc adder4adder43sheet5C34B04AA 1K
R70 adder4adder43sheet5C34B047A adder4adder43sheet5C34B048AorB 10K
R71 adder4adder43sheet5C34B049A adder4adder43sheet5C34B048AorB 10K
Q24 adder4adder43sheet5C34B04AA adder4adder43sheet5C34B048AorB 0 NPN
R75 adder4Vcc adder4adder43sheet5C34B04AB 1K
R73 adder4adder43sheet5C34B049A adder4adder43sheet5C34B049AorB 10K
R74 adder4adder43Cin adder4adder43sheet5C34B049AorB 10K
Q25 adder4adder43sheet5C34B04AB adder4adder43sheet5C34B049AorB 0 NPN
R78 adder4Vcc register4rD3 1K
R76 adder4adder43sheet5C34B04AA adder4adder43sheet5C34B04AAorB 10K
R77 adder4adder43sheet5C34B04AB adder4adder43sheet5C34B04AAorB 10K
Q26 register4rD3 adder4adder43sheet5C34B04AAorB 0 NPN
R81 adder4Vcc adder4adder44Cin 1K
R79 adder4adder43sheet5C34B049A adder4adder43sheet5C34B0CDAorB 10K
R80 adder4adder43sheet5C34B00DA adder4adder43sheet5C34B0CDAorB 10K
Q27 adder4adder44Cin adder4adder43sheet5C34B0CDAorB 0 NPN
R84 adder4Vcc adder4adder44sheet5C34B00DA 1K
R82 adder4A4 adder4adder44sheet5C34AF27AorB 10K
R83 adder4B4 adder4adder44sheet5C34AF27AorB 10K
Q28 adder4adder44sheet5C34B00DA adder4adder44sheet5C34AF27AorB 0 NPN
R87 adder4Vcc adder4adder44sheet5C34B027A 1K
R85 adder4A4 adder4adder44sheet5C34AFF9AorB 10K
R86 adder4adder44sheet5C34B00DA adder4adder44sheet5C34AFF9AorB 10K
Q29 adder4adder44sheet5C34B027A adder4adder44sheet5C34AFF9AorB 0 NPN
R90 adder4Vcc adder4adder44sheet5C34B027B 1K
R88 adder4adder44sheet5C34B00DA adder4adder44sheet5C34B00DAorB 10K
R89 adder4B4 adder4adder44sheet5C34B00DAorB 10K
Q30 adder4adder44sheet5C34B027B adder4adder44sheet5C34B00DAorB 0 NPN
R93 adder4Vcc adder4adder44sheet5C34B047A 1K
R91 adder4adder44sheet5C34B027A adder4adder44sheet5C34B027AorB 10K
R92 adder4adder44sheet5C34B027B adder4adder44sheet5C34B027AorB 10K
Q31 adder4adder44sheet5C34B047A adder4adder44sheet5C34B027AorB 0 NPN
R96 adder4Vcc adder4adder44sheet5C34B049A 1K
R94 adder4adder44sheet5C34B047A adder4adder44sheet5C34B047AorB 10K
R95 adder4adder44Cin adder4adder44sheet5C34B047AorB 10K
Q32 adder4adder44sheet5C34B049A adder4adder44sheet5C34B047AorB 0 NPN
R99 adder4Vcc adder4adder44sheet5C34B04AA 1K
R97 adder4adder44sheet5C34B047A adder4adder44sheet5C34B048AorB 10K
R98 adder4adder44sheet5C34B049A adder4adder44sheet5C34B048AorB 10K
Q33 adder4adder44sheet5C34B04AA adder4adder44sheet5C34B048AorB 0 NPN
R102 adder4Vcc adder4adder44sheet5C34B04AB 1K
R100 adder4adder44sheet5C34B049A adder4adder44sheet5C34B049AorB 10K
R101 adder4adder44Cin adder4adder44sheet5C34B049AorB 10K
Q34 adder4adder44sheet5C34B04AB adder4adder44sheet5C34B049AorB 0 NPN
R105 adder4Vcc register4rD4 1K
R103 adder4adder44sheet5C34B04AA adder4adder44sheet5C34B04AAorB 10K
R104 adder4adder44sheet5C34B04AB adder4adder44sheet5C34B04AAorB 10K
Q35 register4rD4 adder4adder44sheet5C34B04AAorB 0 NPN
R108 adder4Vcc CF 1K
R106 adder4adder44sheet5C34B049A adder4adder44sheet5C34B0CDAorB 10K
R107 adder4adder44sheet5C34B00DA adder4adder44sheet5C34B0CDAorB 10K
Q36 CF adder4adder44sheet5C34B0CDAorB 0 NPN
R111 adder4Vcc adder4A1 1K
R109 register4aregisterflipflop1notd3NQ register4aregisterflipflop1srlatchdsheet5C3630E6AorB 10K
R110 register4aregisterflipflop1NQ register4aregisterflipflop1srlatchdsheet5C3630E6AorB 10K
Q37 adder4A1 register4aregisterflipflop1srlatchdsheet5C3630E6AorB 0 NPN
R114 adder4Vcc register4aregisterflipflop1NQ 1K
R112 adder4A1 register4aregisterflipflop1srlatchdsheet5C3630F6AorB 10K
R113 register4aregisterflipflop1notd2NQ register4aregisterflipflop1srlatchdsheet5C3630F6AorB 10K
Q38 register4aregisterflipflop1NQ register4aregisterflipflop1srlatchdsheet5C3630F6AorB 0 NPN
R116 adder4Vcc register4aregisterflipflop1notd2NQ 1K
R115 register4aregisterflipflop1andd1Q register4aregisterflipflop1notd2Qr 10K
Q39 register4aregisterflipflop1notd2NQ register4aregisterflipflop1notd2Qr 0 NPN
R119 adder4Vcc register4aregisterflipflop1andd1Q 1K
R117 register4aregisterflipflop1andd1sheet5C364DB7A register4aregisterflipflop1andd1sheet5C364DB7AorB 10K
R118 register4aregisterflipflop1andd1sheet5C364DB7B register4aregisterflipflop1andd1sheet5C364DB7AorB 10K
Q40 register4aregisterflipflop1andd1Q register4aregisterflipflop1andd1sheet5C364DB7AorB 0 NPN
R121 adder4Vcc register4aregisterflipflop1andd1sheet5C364DB7A 1K
R120 register4aD1 register4aregisterflipflop1andd1Sheet5C3654CCQr 10K
Q41 register4aregisterflipflop1andd1sheet5C364DB7A register4aregisterflipflop1andd1Sheet5C3654CCQr 0 NPN
R123 adder4Vcc register4aregisterflipflop1andd1sheet5C364DB7B 1K
R122 register4aCLK register4aregisterflipflop1andd1sheet5C366192Qr 10K
Q42 register4aregisterflipflop1andd1sheet5C364DB7B register4aregisterflipflop1andd1sheet5C366192Qr 0 NPN
R125 adder4Vcc register4aregisterflipflop1andd2B 1K
R124 register4aD1 register4aregisterflipflop1notd1Qr 10K
Q43 register4aregisterflipflop1andd2B register4aregisterflipflop1notd1Qr 0 NPN
R127 adder4Vcc register4aregisterflipflop1notd3NQ 1K
R126 register4aregisterflipflop1andd2Q register4aregisterflipflop1notd3Qr 10K
Q44 register4aregisterflipflop1notd3NQ register4aregisterflipflop1notd3Qr 0 NPN
R130 adder4Vcc register4aregisterflipflop1andd2Q 1K
R128 register4aregisterflipflop1andd2sheet5C364DB7A register4aregisterflipflop1andd2sheet5C364DB7AorB 10K
R129 register4aregisterflipflop1andd2sheet5C364DB7B register4aregisterflipflop1andd2sheet5C364DB7AorB 10K
Q45 register4aregisterflipflop1andd2Q register4aregisterflipflop1andd2sheet5C364DB7AorB 0 NPN
R132 adder4Vcc register4aregisterflipflop1andd2sheet5C364DB7A 1K
R131 register4aCLK register4aregisterflipflop1andd2Sheet5C3654CCQr 10K
Q46 register4aregisterflipflop1andd2sheet5C364DB7A register4aregisterflipflop1andd2Sheet5C3654CCQr 0 NPN
R134 adder4Vcc register4aregisterflipflop1andd2sheet5C364DB7B 1K
R133 register4aregisterflipflop1andd2B register4aregisterflipflop1andd2sheet5C366192Qr 10K
Q47 register4aregisterflipflop1andd2sheet5C364DB7B register4aregisterflipflop1andd2sheet5C366192Qr 0 NPN
R137 adder4Vcc adder4A2 1K
R135 register4aregisterflipflop2notd3NQ register4aregisterflipflop2srlatchdsheet5C3630E6AorB 10K
R136 register4aregisterflipflop2NQ register4aregisterflipflop2srlatchdsheet5C3630E6AorB 10K
Q48 adder4A2 register4aregisterflipflop2srlatchdsheet5C3630E6AorB 0 NPN
R140 adder4Vcc register4aregisterflipflop2NQ 1K
R138 adder4A2 register4aregisterflipflop2srlatchdsheet5C3630F6AorB 10K
R139 register4aregisterflipflop2notd2NQ register4aregisterflipflop2srlatchdsheet5C3630F6AorB 10K
Q49 register4aregisterflipflop2NQ register4aregisterflipflop2srlatchdsheet5C3630F6AorB 0 NPN
R142 adder4Vcc register4aregisterflipflop2notd2NQ 1K
R141 register4aregisterflipflop2andd1Q register4aregisterflipflop2notd2Qr 10K
Q50 register4aregisterflipflop2notd2NQ register4aregisterflipflop2notd2Qr 0 NPN
R145 adder4Vcc register4aregisterflipflop2andd1Q 1K
R143 register4aregisterflipflop2andd1sheet5C364DB7A register4aregisterflipflop2andd1sheet5C364DB7AorB 10K
R144 register4aregisterflipflop2andd1sheet5C364DB7B register4aregisterflipflop2andd1sheet5C364DB7AorB 10K
Q51 register4aregisterflipflop2andd1Q register4aregisterflipflop2andd1sheet5C364DB7AorB 0 NPN
R147 adder4Vcc register4aregisterflipflop2andd1sheet5C364DB7A 1K
R146 register4aD2 register4aregisterflipflop2andd1Sheet5C3654CCQr 10K
Q52 register4aregisterflipflop2andd1sheet5C364DB7A register4aregisterflipflop2andd1Sheet5C3654CCQr 0 NPN
R149 adder4Vcc register4aregisterflipflop2andd1sheet5C364DB7B 1K
R148 register4aCLK register4aregisterflipflop2andd1sheet5C366192Qr 10K
Q53 register4aregisterflipflop2andd1sheet5C364DB7B register4aregisterflipflop2andd1sheet5C366192Qr 0 NPN
R151 adder4Vcc register4aregisterflipflop2andd2B 1K
R150 register4aD2 register4aregisterflipflop2notd1Qr 10K
Q54 register4aregisterflipflop2andd2B register4aregisterflipflop2notd1Qr 0 NPN
R153 adder4Vcc register4aregisterflipflop2notd3NQ 1K
R152 register4aregisterflipflop2andd2Q register4aregisterflipflop2notd3Qr 10K
Q55 register4aregisterflipflop2notd3NQ register4aregisterflipflop2notd3Qr 0 NPN
R156 adder4Vcc register4aregisterflipflop2andd2Q 1K
R154 register4aregisterflipflop2andd2sheet5C364DB7A register4aregisterflipflop2andd2sheet5C364DB7AorB 10K
R155 register4aregisterflipflop2andd2sheet5C364DB7B register4aregisterflipflop2andd2sheet5C364DB7AorB 10K
Q56 register4aregisterflipflop2andd2Q register4aregisterflipflop2andd2sheet5C364DB7AorB 0 NPN
R158 adder4Vcc register4aregisterflipflop2andd2sheet5C364DB7A 1K
R157 register4aCLK register4aregisterflipflop2andd2Sheet5C3654CCQr 10K
Q57 register4aregisterflipflop2andd2sheet5C364DB7A register4aregisterflipflop2andd2Sheet5C3654CCQr 0 NPN
R160 adder4Vcc register4aregisterflipflop2andd2sheet5C364DB7B 1K
R159 register4aregisterflipflop2andd2B register4aregisterflipflop2andd2sheet5C366192Qr 10K
Q58 register4aregisterflipflop2andd2sheet5C364DB7B register4aregisterflipflop2andd2sheet5C366192Qr 0 NPN
R163 adder4Vcc adder4A3 1K
R161 register4aregisterflipflop3notd3NQ register4aregisterflipflop3srlatchdsheet5C3630E6AorB 10K
R162 register4aregisterflipflop3NQ register4aregisterflipflop3srlatchdsheet5C3630E6AorB 10K
Q59 adder4A3 register4aregisterflipflop3srlatchdsheet5C3630E6AorB 0 NPN
R166 adder4Vcc register4aregisterflipflop3NQ 1K
R164 adder4A3 register4aregisterflipflop3srlatchdsheet5C3630F6AorB 10K
R165 register4aregisterflipflop3notd2NQ register4aregisterflipflop3srlatchdsheet5C3630F6AorB 10K
Q60 register4aregisterflipflop3NQ register4aregisterflipflop3srlatchdsheet5C3630F6AorB 0 NPN
R168 adder4Vcc register4aregisterflipflop3notd2NQ 1K
R167 register4aregisterflipflop3andd1Q register4aregisterflipflop3notd2Qr 10K
Q61 register4aregisterflipflop3notd2NQ register4aregisterflipflop3notd2Qr 0 NPN
R171 adder4Vcc register4aregisterflipflop3andd1Q 1K
R169 register4aregisterflipflop3andd1sheet5C364DB7A register4aregisterflipflop3andd1sheet5C364DB7AorB 10K
R170 register4aregisterflipflop3andd1sheet5C364DB7B register4aregisterflipflop3andd1sheet5C364DB7AorB 10K
Q62 register4aregisterflipflop3andd1Q register4aregisterflipflop3andd1sheet5C364DB7AorB 0 NPN
R173 adder4Vcc register4aregisterflipflop3andd1sheet5C364DB7A 1K
R172 register4aD3 register4aregisterflipflop3andd1Sheet5C3654CCQr 10K
Q63 register4aregisterflipflop3andd1sheet5C364DB7A register4aregisterflipflop3andd1Sheet5C3654CCQr 0 NPN
R175 adder4Vcc register4aregisterflipflop3andd1sheet5C364DB7B 1K
R174 register4aCLK register4aregisterflipflop3andd1sheet5C366192Qr 10K
Q64 register4aregisterflipflop3andd1sheet5C364DB7B register4aregisterflipflop3andd1sheet5C366192Qr 0 NPN
R177 adder4Vcc register4aregisterflipflop3andd2B 1K
R176 register4aD3 register4aregisterflipflop3notd1Qr 10K
Q65 register4aregisterflipflop3andd2B register4aregisterflipflop3notd1Qr 0 NPN
R179 adder4Vcc register4aregisterflipflop3notd3NQ 1K
R178 register4aregisterflipflop3andd2Q register4aregisterflipflop3notd3Qr 10K
Q66 register4aregisterflipflop3notd3NQ register4aregisterflipflop3notd3Qr 0 NPN
R182 adder4Vcc register4aregisterflipflop3andd2Q 1K
R180 register4aregisterflipflop3andd2sheet5C364DB7A register4aregisterflipflop3andd2sheet5C364DB7AorB 10K
R181 register4aregisterflipflop3andd2sheet5C364DB7B register4aregisterflipflop3andd2sheet5C364DB7AorB 10K
Q67 register4aregisterflipflop3andd2Q register4aregisterflipflop3andd2sheet5C364DB7AorB 0 NPN
R184 adder4Vcc register4aregisterflipflop3andd2sheet5C364DB7A 1K
R183 register4aCLK register4aregisterflipflop3andd2Sheet5C3654CCQr 10K
Q68 register4aregisterflipflop3andd2sheet5C364DB7A register4aregisterflipflop3andd2Sheet5C3654CCQr 0 NPN
R186 adder4Vcc register4aregisterflipflop3andd2sheet5C364DB7B 1K
R185 register4aregisterflipflop3andd2B register4aregisterflipflop3andd2sheet5C366192Qr 10K
Q69 register4aregisterflipflop3andd2sheet5C364DB7B register4aregisterflipflop3andd2sheet5C366192Qr 0 NPN
R189 adder4Vcc adder4A4 1K
R187 register4aregisterflipflop4notd3NQ register4aregisterflipflop4srlatchdsheet5C3630E6AorB 10K
R188 register4aregisterflipflop4NQ register4aregisterflipflop4srlatchdsheet5C3630E6AorB 10K
Q70 adder4A4 register4aregisterflipflop4srlatchdsheet5C3630E6AorB 0 NPN
R192 adder4Vcc register4aregisterflipflop4NQ 1K
R190 adder4A4 register4aregisterflipflop4srlatchdsheet5C3630F6AorB 10K
R191 register4aregisterflipflop4notd2NQ register4aregisterflipflop4srlatchdsheet5C3630F6AorB 10K
Q71 register4aregisterflipflop4NQ register4aregisterflipflop4srlatchdsheet5C3630F6AorB 0 NPN
R194 adder4Vcc register4aregisterflipflop4notd2NQ 1K
R193 register4aregisterflipflop4andd1Q register4aregisterflipflop4notd2Qr 10K
Q72 register4aregisterflipflop4notd2NQ register4aregisterflipflop4notd2Qr 0 NPN
R197 adder4Vcc register4aregisterflipflop4andd1Q 1K
R195 register4aregisterflipflop4andd1sheet5C364DB7A register4aregisterflipflop4andd1sheet5C364DB7AorB 10K
R196 register4aregisterflipflop4andd1sheet5C364DB7B register4aregisterflipflop4andd1sheet5C364DB7AorB 10K
Q73 register4aregisterflipflop4andd1Q register4aregisterflipflop4andd1sheet5C364DB7AorB 0 NPN
R199 adder4Vcc register4aregisterflipflop4andd1sheet5C364DB7A 1K
R198 register4aD4 register4aregisterflipflop4andd1Sheet5C3654CCQr 10K
Q74 register4aregisterflipflop4andd1sheet5C364DB7A register4aregisterflipflop4andd1Sheet5C3654CCQr 0 NPN
R201 adder4Vcc register4aregisterflipflop4andd1sheet5C364DB7B 1K
R200 register4aCLK register4aregisterflipflop4andd1sheet5C366192Qr 10K
Q75 register4aregisterflipflop4andd1sheet5C364DB7B register4aregisterflipflop4andd1sheet5C366192Qr 0 NPN
R203 adder4Vcc register4aregisterflipflop4andd2B 1K
R202 register4aD4 register4aregisterflipflop4notd1Qr 10K
Q76 register4aregisterflipflop4andd2B register4aregisterflipflop4notd1Qr 0 NPN
R205 adder4Vcc register4aregisterflipflop4notd3NQ 1K
R204 register4aregisterflipflop4andd2Q register4aregisterflipflop4notd3Qr 10K
Q77 register4aregisterflipflop4notd3NQ register4aregisterflipflop4notd3Qr 0 NPN
R208 adder4Vcc register4aregisterflipflop4andd2Q 1K
R206 register4aregisterflipflop4andd2sheet5C364DB7A register4aregisterflipflop4andd2sheet5C364DB7AorB 10K
R207 register4aregisterflipflop4andd2sheet5C364DB7B register4aregisterflipflop4andd2sheet5C364DB7AorB 10K
Q78 register4aregisterflipflop4andd2Q register4aregisterflipflop4andd2sheet5C364DB7AorB 0 NPN
R210 adder4Vcc register4aregisterflipflop4andd2sheet5C364DB7A 1K
R209 register4aCLK register4aregisterflipflop4andd2Sheet5C3654CCQr 10K
Q79 register4aregisterflipflop4andd2sheet5C364DB7A register4aregisterflipflop4andd2Sheet5C3654CCQr 0 NPN
R212 adder4Vcc register4aregisterflipflop4andd2sheet5C364DB7B 1K
R211 register4aregisterflipflop4andd2B register4aregisterflipflop4andd2sheet5C366192Qr 10K
Q80 register4aregisterflipflop4andd2sheet5C364DB7B register4aregisterflipflop4andd2sheet5C366192Qr 0 NPN
R215 adder4Vcc adder4B1 1K
R213 register4bregisterflipflop1notd3NQ register4bregisterflipflop1srlatchdsheet5C3630E6AorB 10K
R214 register4bregisterflipflop1NQ register4bregisterflipflop1srlatchdsheet5C3630E6AorB 10K
Q81 adder4B1 register4bregisterflipflop1srlatchdsheet5C3630E6AorB 0 NPN
R218 adder4Vcc register4bregisterflipflop1NQ 1K
R216 adder4B1 register4bregisterflipflop1srlatchdsheet5C3630F6AorB 10K
R217 register4bregisterflipflop1notd2NQ register4bregisterflipflop1srlatchdsheet5C3630F6AorB 10K
Q82 register4bregisterflipflop1NQ register4bregisterflipflop1srlatchdsheet5C3630F6AorB 0 NPN
R220 adder4Vcc register4bregisterflipflop1notd2NQ 1K
R219 register4bregisterflipflop1andd1Q register4bregisterflipflop1notd2Qr 10K
Q83 register4bregisterflipflop1notd2NQ register4bregisterflipflop1notd2Qr 0 NPN
R223 adder4Vcc register4bregisterflipflop1andd1Q 1K
R221 register4bregisterflipflop1andd1sheet5C364DB7A register4bregisterflipflop1andd1sheet5C364DB7AorB 10K
R222 register4bregisterflipflop1andd1sheet5C364DB7B register4bregisterflipflop1andd1sheet5C364DB7AorB 10K
Q84 register4bregisterflipflop1andd1Q register4bregisterflipflop1andd1sheet5C364DB7AorB 0 NPN
R225 adder4Vcc register4bregisterflipflop1andd1sheet5C364DB7A 1K
R224 register4bD1 register4bregisterflipflop1andd1Sheet5C3654CCQr 10K
Q85 register4bregisterflipflop1andd1sheet5C364DB7A register4bregisterflipflop1andd1Sheet5C3654CCQr 0 NPN
R227 adder4Vcc register4bregisterflipflop1andd1sheet5C364DB7B 1K
R226 register4aCLK register4bregisterflipflop1andd1sheet5C366192Qr 10K
Q86 register4bregisterflipflop1andd1sheet5C364DB7B register4bregisterflipflop1andd1sheet5C366192Qr 0 NPN
R229 adder4Vcc register4bregisterflipflop1andd2B 1K
R228 register4bD1 register4bregisterflipflop1notd1Qr 10K
Q87 register4bregisterflipflop1andd2B register4bregisterflipflop1notd1Qr 0 NPN
R231 adder4Vcc register4bregisterflipflop1notd3NQ 1K
R230 register4bregisterflipflop1andd2Q register4bregisterflipflop1notd3Qr 10K
Q88 register4bregisterflipflop1notd3NQ register4bregisterflipflop1notd3Qr 0 NPN
R234 adder4Vcc register4bregisterflipflop1andd2Q 1K
R232 register4bregisterflipflop1andd2sheet5C364DB7A register4bregisterflipflop1andd2sheet5C364DB7AorB 10K
R233 register4bregisterflipflop1andd2sheet5C364DB7B register4bregisterflipflop1andd2sheet5C364DB7AorB 10K
Q89 register4bregisterflipflop1andd2Q register4bregisterflipflop1andd2sheet5C364DB7AorB 0 NPN
R236 adder4Vcc register4bregisterflipflop1andd2sheet5C364DB7A 1K
R235 register4aCLK register4bregisterflipflop1andd2Sheet5C3654CCQr 10K
Q90 register4bregisterflipflop1andd2sheet5C364DB7A register4bregisterflipflop1andd2Sheet5C3654CCQr 0 NPN
R238 adder4Vcc register4bregisterflipflop1andd2sheet5C364DB7B 1K
R237 register4bregisterflipflop1andd2B register4bregisterflipflop1andd2sheet5C366192Qr 10K
Q91 register4bregisterflipflop1andd2sheet5C364DB7B register4bregisterflipflop1andd2sheet5C366192Qr 0 NPN
R241 adder4Vcc adder4B2 1K
R239 register4bregisterflipflop2notd3NQ register4bregisterflipflop2srlatchdsheet5C3630E6AorB 10K
R240 register4bregisterflipflop2NQ register4bregisterflipflop2srlatchdsheet5C3630E6AorB 10K
Q92 adder4B2 register4bregisterflipflop2srlatchdsheet5C3630E6AorB 0 NPN
R244 adder4Vcc register4bregisterflipflop2NQ 1K
R242 adder4B2 register4bregisterflipflop2srlatchdsheet5C3630F6AorB 10K
R243 register4bregisterflipflop2notd2NQ register4bregisterflipflop2srlatchdsheet5C3630F6AorB 10K
Q93 register4bregisterflipflop2NQ register4bregisterflipflop2srlatchdsheet5C3630F6AorB 0 NPN
R246 adder4Vcc register4bregisterflipflop2notd2NQ 1K
R245 register4bregisterflipflop2andd1Q register4bregisterflipflop2notd2Qr 10K
Q94 register4bregisterflipflop2notd2NQ register4bregisterflipflop2notd2Qr 0 NPN
R249 adder4Vcc register4bregisterflipflop2andd1Q 1K
R247 register4bregisterflipflop2andd1sheet5C364DB7A register4bregisterflipflop2andd1sheet5C364DB7AorB 10K
R248 register4bregisterflipflop2andd1sheet5C364DB7B register4bregisterflipflop2andd1sheet5C364DB7AorB 10K
Q95 register4bregisterflipflop2andd1Q register4bregisterflipflop2andd1sheet5C364DB7AorB 0 NPN
R251 adder4Vcc register4bregisterflipflop2andd1sheet5C364DB7A 1K
R250 register4bD2 register4bregisterflipflop2andd1Sheet5C3654CCQr 10K
Q96 register4bregisterflipflop2andd1sheet5C364DB7A register4bregisterflipflop2andd1Sheet5C3654CCQr 0 NPN
R253 adder4Vcc register4bregisterflipflop2andd1sheet5C364DB7B 1K
R252 register4aCLK register4bregisterflipflop2andd1sheet5C366192Qr 10K
Q97 register4bregisterflipflop2andd1sheet5C364DB7B register4bregisterflipflop2andd1sheet5C366192Qr 0 NPN
R255 adder4Vcc register4bregisterflipflop2andd2B 1K
R254 register4bD2 register4bregisterflipflop2notd1Qr 10K
Q98 register4bregisterflipflop2andd2B register4bregisterflipflop2notd1Qr 0 NPN
R257 adder4Vcc register4bregisterflipflop2notd3NQ 1K
R256 register4bregisterflipflop2andd2Q register4bregisterflipflop2notd3Qr 10K
Q99 register4bregisterflipflop2notd3NQ register4bregisterflipflop2notd3Qr 0 NPN
R260 adder4Vcc register4bregisterflipflop2andd2Q 1K
R258 register4bregisterflipflop2andd2sheet5C364DB7A register4bregisterflipflop2andd2sheet5C364DB7AorB 10K
R259 register4bregisterflipflop2andd2sheet5C364DB7B register4bregisterflipflop2andd2sheet5C364DB7AorB 10K
Q100 register4bregisterflipflop2andd2Q register4bregisterflipflop2andd2sheet5C364DB7AorB 0 NPN
R262 adder4Vcc register4bregisterflipflop2andd2sheet5C364DB7A 1K
R261 register4aCLK register4bregisterflipflop2andd2Sheet5C3654CCQr 10K
Q101 register4bregisterflipflop2andd2sheet5C364DB7A register4bregisterflipflop2andd2Sheet5C3654CCQr 0 NPN
R264 adder4Vcc register4bregisterflipflop2andd2sheet5C364DB7B 1K
R263 register4bregisterflipflop2andd2B register4bregisterflipflop2andd2sheet5C366192Qr 10K
Q102 register4bregisterflipflop2andd2sheet5C364DB7B register4bregisterflipflop2andd2sheet5C366192Qr 0 NPN
R267 adder4Vcc adder4B3 1K
R265 register4bregisterflipflop3notd3NQ register4bregisterflipflop3srlatchdsheet5C3630E6AorB 10K
R266 register4bregisterflipflop3NQ register4bregisterflipflop3srlatchdsheet5C3630E6AorB 10K
Q103 adder4B3 register4bregisterflipflop3srlatchdsheet5C3630E6AorB 0 NPN
R270 adder4Vcc register4bregisterflipflop3NQ 1K
R268 adder4B3 register4bregisterflipflop3srlatchdsheet5C3630F6AorB 10K
R269 register4bregisterflipflop3notd2NQ register4bregisterflipflop3srlatchdsheet5C3630F6AorB 10K
Q104 register4bregisterflipflop3NQ register4bregisterflipflop3srlatchdsheet5C3630F6AorB 0 NPN
R272 adder4Vcc register4bregisterflipflop3notd2NQ 1K
R271 register4bregisterflipflop3andd1Q register4bregisterflipflop3notd2Qr 10K
Q105 register4bregisterflipflop3notd2NQ register4bregisterflipflop3notd2Qr 0 NPN
R275 adder4Vcc register4bregisterflipflop3andd1Q 1K
R273 register4bregisterflipflop3andd1sheet5C364DB7A register4bregisterflipflop3andd1sheet5C364DB7AorB 10K
R274 register4bregisterflipflop3andd1sheet5C364DB7B register4bregisterflipflop3andd1sheet5C364DB7AorB 10K
Q106 register4bregisterflipflop3andd1Q register4bregisterflipflop3andd1sheet5C364DB7AorB 0 NPN
R277 adder4Vcc register4bregisterflipflop3andd1sheet5C364DB7A 1K
R276 register4bD3 register4bregisterflipflop3andd1Sheet5C3654CCQr 10K
Q107 register4bregisterflipflop3andd1sheet5C364DB7A register4bregisterflipflop3andd1Sheet5C3654CCQr 0 NPN
R279 adder4Vcc register4bregisterflipflop3andd1sheet5C364DB7B 1K
R278 register4aCLK register4bregisterflipflop3andd1sheet5C366192Qr 10K
Q108 register4bregisterflipflop3andd1sheet5C364DB7B register4bregisterflipflop3andd1sheet5C366192Qr 0 NPN
R281 adder4Vcc register4bregisterflipflop3andd2B 1K
R280 register4bD3 register4bregisterflipflop3notd1Qr 10K
Q109 register4bregisterflipflop3andd2B register4bregisterflipflop3notd1Qr 0 NPN
R283 adder4Vcc register4bregisterflipflop3notd3NQ 1K
R282 register4bregisterflipflop3andd2Q register4bregisterflipflop3notd3Qr 10K
Q110 register4bregisterflipflop3notd3NQ register4bregisterflipflop3notd3Qr 0 NPN
R286 adder4Vcc register4bregisterflipflop3andd2Q 1K
R284 register4bregisterflipflop3andd2sheet5C364DB7A register4bregisterflipflop3andd2sheet5C364DB7AorB 10K
R285 register4bregisterflipflop3andd2sheet5C364DB7B register4bregisterflipflop3andd2sheet5C364DB7AorB 10K
Q111 register4bregisterflipflop3andd2Q register4bregisterflipflop3andd2sheet5C364DB7AorB 0 NPN
R288 adder4Vcc register4bregisterflipflop3andd2sheet5C364DB7A 1K
R287 register4aCLK register4bregisterflipflop3andd2Sheet5C3654CCQr 10K
Q112 register4bregisterflipflop3andd2sheet5C364DB7A register4bregisterflipflop3andd2Sheet5C3654CCQr 0 NPN
R290 adder4Vcc register4bregisterflipflop3andd2sheet5C364DB7B 1K
R289 register4bregisterflipflop3andd2B register4bregisterflipflop3andd2sheet5C366192Qr 10K
Q113 register4bregisterflipflop3andd2sheet5C364DB7B register4bregisterflipflop3andd2sheet5C366192Qr 0 NPN
R293 adder4Vcc adder4B4 1K
R291 register4bregisterflipflop4notd3NQ register4bregisterflipflop4srlatchdsheet5C3630E6AorB 10K
R292 register4bregisterflipflop4NQ register4bregisterflipflop4srlatchdsheet5C3630E6AorB 10K
Q114 adder4B4 register4bregisterflipflop4srlatchdsheet5C3630E6AorB 0 NPN
R296 adder4Vcc register4bregisterflipflop4NQ 1K
R294 adder4B4 register4bregisterflipflop4srlatchdsheet5C3630F6AorB 10K
R295 register4bregisterflipflop4notd2NQ register4bregisterflipflop4srlatchdsheet5C3630F6AorB 10K
Q115 register4bregisterflipflop4NQ register4bregisterflipflop4srlatchdsheet5C3630F6AorB 0 NPN
R298 adder4Vcc register4bregisterflipflop4notd2NQ 1K
R297 register4bregisterflipflop4andd1Q register4bregisterflipflop4notd2Qr 10K
Q116 register4bregisterflipflop4notd2NQ register4bregisterflipflop4notd2Qr 0 NPN
R301 adder4Vcc register4bregisterflipflop4andd1Q 1K
R299 register4bregisterflipflop4andd1sheet5C364DB7A register4bregisterflipflop4andd1sheet5C364DB7AorB 10K
R300 register4bregisterflipflop4andd1sheet5C364DB7B register4bregisterflipflop4andd1sheet5C364DB7AorB 10K
Q117 register4bregisterflipflop4andd1Q register4bregisterflipflop4andd1sheet5C364DB7AorB 0 NPN
R303 adder4Vcc register4bregisterflipflop4andd1sheet5C364DB7A 1K
R302 register4bD4 register4bregisterflipflop4andd1Sheet5C3654CCQr 10K
Q118 register4bregisterflipflop4andd1sheet5C364DB7A register4bregisterflipflop4andd1Sheet5C3654CCQr 0 NPN
R305 adder4Vcc register4bregisterflipflop4andd1sheet5C364DB7B 1K
R304 register4aCLK register4bregisterflipflop4andd1sheet5C366192Qr 10K
Q119 register4bregisterflipflop4andd1sheet5C364DB7B register4bregisterflipflop4andd1sheet5C366192Qr 0 NPN
R307 adder4Vcc register4bregisterflipflop4andd2B 1K
R306 register4bD4 register4bregisterflipflop4notd1Qr 10K
Q120 register4bregisterflipflop4andd2B register4bregisterflipflop4notd1Qr 0 NPN
R309 adder4Vcc register4bregisterflipflop4notd3NQ 1K
R308 register4bregisterflipflop4andd2Q register4bregisterflipflop4notd3Qr 10K
Q121 register4bregisterflipflop4notd3NQ register4bregisterflipflop4notd3Qr 0 NPN
R312 adder4Vcc register4bregisterflipflop4andd2Q 1K
R310 register4bregisterflipflop4andd2sheet5C364DB7A register4bregisterflipflop4andd2sheet5C364DB7AorB 10K
R311 register4bregisterflipflop4andd2sheet5C364DB7B register4bregisterflipflop4andd2sheet5C364DB7AorB 10K
Q122 register4bregisterflipflop4andd2Q register4bregisterflipflop4andd2sheet5C364DB7AorB 0 NPN
R314 adder4Vcc register4bregisterflipflop4andd2sheet5C364DB7A 1K
R313 register4aCLK register4bregisterflipflop4andd2Sheet5C3654CCQr 10K
Q123 register4bregisterflipflop4andd2sheet5C364DB7A register4bregisterflipflop4andd2Sheet5C3654CCQr 0 NPN
R316 adder4Vcc register4bregisterflipflop4andd2sheet5C364DB7B 1K
R315 register4bregisterflipflop4andd2B register4bregisterflipflop4andd2sheet5C366192Qr 10K
Q124 register4bregisterflipflop4andd2sheet5C364DB7B register4bregisterflipflop4andd2sheet5C366192Qr 0 NPN
R319 adder4Vcc register4rQ1 1K
R317 register4rregisterflipflop1notd3NQ register4rregisterflipflop1srlatchdsheet5C3630E6AorB 10K
R318 register4rregisterflipflop1NQ register4rregisterflipflop1srlatchdsheet5C3630E6AorB 10K
Q125 register4rQ1 register4rregisterflipflop1srlatchdsheet5C3630E6AorB 0 NPN
R322 adder4Vcc register4rregisterflipflop1NQ 1K
R320 register4rQ1 register4rregisterflipflop1srlatchdsheet5C3630F6AorB 10K
R321 register4rregisterflipflop1notd2NQ register4rregisterflipflop1srlatchdsheet5C3630F6AorB 10K
Q126 register4rregisterflipflop1NQ register4rregisterflipflop1srlatchdsheet5C3630F6AorB 0 NPN
R324 adder4Vcc register4rregisterflipflop1notd2NQ 1K
R323 register4rregisterflipflop1andd1Q register4rregisterflipflop1notd2Qr 10K
Q127 register4rregisterflipflop1notd2NQ register4rregisterflipflop1notd2Qr 0 NPN
R327 adder4Vcc register4rregisterflipflop1andd1Q 1K
R325 register4rregisterflipflop1andd1sheet5C364DB7A register4rregisterflipflop1andd1sheet5C364DB7AorB 10K
R326 register4rregisterflipflop1andd1sheet5C364DB7B register4rregisterflipflop1andd1sheet5C364DB7AorB 10K
Q128 register4rregisterflipflop1andd1Q register4rregisterflipflop1andd1sheet5C364DB7AorB 0 NPN
R329 adder4Vcc register4rregisterflipflop1andd1sheet5C364DB7A 1K
R328 register4rD1 register4rregisterflipflop1andd1Sheet5C3654CCQr 10K
Q129 register4rregisterflipflop1andd1sheet5C364DB7A register4rregisterflipflop1andd1Sheet5C3654CCQr 0 NPN
R331 adder4Vcc register4rregisterflipflop1andd1sheet5C364DB7B 1K
R330 register4aCLK register4rregisterflipflop1andd1sheet5C366192Qr 10K
Q130 register4rregisterflipflop1andd1sheet5C364DB7B register4rregisterflipflop1andd1sheet5C366192Qr 0 NPN
R333 adder4Vcc register4rregisterflipflop1andd2B 1K
R332 register4rD1 register4rregisterflipflop1notd1Qr 10K
Q131 register4rregisterflipflop1andd2B register4rregisterflipflop1notd1Qr 0 NPN
R335 adder4Vcc register4rregisterflipflop1notd3NQ 1K
R334 register4rregisterflipflop1andd2Q register4rregisterflipflop1notd3Qr 10K
Q132 register4rregisterflipflop1notd3NQ register4rregisterflipflop1notd3Qr 0 NPN
R338 adder4Vcc register4rregisterflipflop1andd2Q 1K
R336 register4rregisterflipflop1andd2sheet5C364DB7A register4rregisterflipflop1andd2sheet5C364DB7AorB 10K
R337 register4rregisterflipflop1andd2sheet5C364DB7B register4rregisterflipflop1andd2sheet5C364DB7AorB 10K
Q133 register4rregisterflipflop1andd2Q register4rregisterflipflop1andd2sheet5C364DB7AorB 0 NPN
R340 adder4Vcc register4rregisterflipflop1andd2sheet5C364DB7A 1K
R339 register4aCLK register4rregisterflipflop1andd2Sheet5C3654CCQr 10K
Q134 register4rregisterflipflop1andd2sheet5C364DB7A register4rregisterflipflop1andd2Sheet5C3654CCQr 0 NPN
R342 adder4Vcc register4rregisterflipflop1andd2sheet5C364DB7B 1K
R341 register4rregisterflipflop1andd2B register4rregisterflipflop1andd2sheet5C366192Qr 10K
Q135 register4rregisterflipflop1andd2sheet5C364DB7B register4rregisterflipflop1andd2sheet5C366192Qr 0 NPN
R345 adder4Vcc register4rQ2 1K
R343 register4rregisterflipflop2notd3NQ register4rregisterflipflop2srlatchdsheet5C3630E6AorB 10K
R344 register4rregisterflipflop2NQ register4rregisterflipflop2srlatchdsheet5C3630E6AorB 10K
Q136 register4rQ2 register4rregisterflipflop2srlatchdsheet5C3630E6AorB 0 NPN
R348 adder4Vcc register4rregisterflipflop2NQ 1K
R346 register4rQ2 register4rregisterflipflop2srlatchdsheet5C3630F6AorB 10K
R347 register4rregisterflipflop2notd2NQ register4rregisterflipflop2srlatchdsheet5C3630F6AorB 10K
Q137 register4rregisterflipflop2NQ register4rregisterflipflop2srlatchdsheet5C3630F6AorB 0 NPN
R350 adder4Vcc register4rregisterflipflop2notd2NQ 1K
R349 register4rregisterflipflop2andd1Q register4rregisterflipflop2notd2Qr 10K
Q138 register4rregisterflipflop2notd2NQ register4rregisterflipflop2notd2Qr 0 NPN
R353 adder4Vcc register4rregisterflipflop2andd1Q 1K
R351 register4rregisterflipflop2andd1sheet5C364DB7A register4rregisterflipflop2andd1sheet5C364DB7AorB 10K
R352 register4rregisterflipflop2andd1sheet5C364DB7B register4rregisterflipflop2andd1sheet5C364DB7AorB 10K
Q139 register4rregisterflipflop2andd1Q register4rregisterflipflop2andd1sheet5C364DB7AorB 0 NPN
R355 adder4Vcc register4rregisterflipflop2andd1sheet5C364DB7A 1K
R354 register4rD2 register4rregisterflipflop2andd1Sheet5C3654CCQr 10K
Q140 register4rregisterflipflop2andd1sheet5C364DB7A register4rregisterflipflop2andd1Sheet5C3654CCQr 0 NPN
R357 adder4Vcc register4rregisterflipflop2andd1sheet5C364DB7B 1K
R356 register4aCLK register4rregisterflipflop2andd1sheet5C366192Qr 10K
Q141 register4rregisterflipflop2andd1sheet5C364DB7B register4rregisterflipflop2andd1sheet5C366192Qr 0 NPN
R359 adder4Vcc register4rregisterflipflop2andd2B 1K
R358 register4rD2 register4rregisterflipflop2notd1Qr 10K
Q142 register4rregisterflipflop2andd2B register4rregisterflipflop2notd1Qr 0 NPN
R361 adder4Vcc register4rregisterflipflop2notd3NQ 1K
R360 register4rregisterflipflop2andd2Q register4rregisterflipflop2notd3Qr 10K
Q143 register4rregisterflipflop2notd3NQ register4rregisterflipflop2notd3Qr 0 NPN
R364 adder4Vcc register4rregisterflipflop2andd2Q 1K
R362 register4rregisterflipflop2andd2sheet5C364DB7A register4rregisterflipflop2andd2sheet5C364DB7AorB 10K
R363 register4rregisterflipflop2andd2sheet5C364DB7B register4rregisterflipflop2andd2sheet5C364DB7AorB 10K
Q144 register4rregisterflipflop2andd2Q register4rregisterflipflop2andd2sheet5C364DB7AorB 0 NPN
R366 adder4Vcc register4rregisterflipflop2andd2sheet5C364DB7A 1K
R365 register4aCLK register4rregisterflipflop2andd2Sheet5C3654CCQr 10K
Q145 register4rregisterflipflop2andd2sheet5C364DB7A register4rregisterflipflop2andd2Sheet5C3654CCQr 0 NPN
R368 adder4Vcc register4rregisterflipflop2andd2sheet5C364DB7B 1K
R367 register4rregisterflipflop2andd2B register4rregisterflipflop2andd2sheet5C366192Qr 10K
Q146 register4rregisterflipflop2andd2sheet5C364DB7B register4rregisterflipflop2andd2sheet5C366192Qr 0 NPN
R371 adder4Vcc register4rQ3 1K
R369 register4rregisterflipflop3notd3NQ register4rregisterflipflop3srlatchdsheet5C3630E6AorB 10K
R370 register4rregisterflipflop3NQ register4rregisterflipflop3srlatchdsheet5C3630E6AorB 10K
Q147 register4rQ3 register4rregisterflipflop3srlatchdsheet5C3630E6AorB 0 NPN
R374 adder4Vcc register4rregisterflipflop3NQ 1K
R372 register4rQ3 register4rregisterflipflop3srlatchdsheet5C3630F6AorB 10K
R373 register4rregisterflipflop3notd2NQ register4rregisterflipflop3srlatchdsheet5C3630F6AorB 10K
Q148 register4rregisterflipflop3NQ register4rregisterflipflop3srlatchdsheet5C3630F6AorB 0 NPN
R376 adder4Vcc register4rregisterflipflop3notd2NQ 1K
R375 register4rregisterflipflop3andd1Q register4rregisterflipflop3notd2Qr 10K
Q149 register4rregisterflipflop3notd2NQ register4rregisterflipflop3notd2Qr 0 NPN
R379 adder4Vcc register4rregisterflipflop3andd1Q 1K
R377 register4rregisterflipflop3andd1sheet5C364DB7A register4rregisterflipflop3andd1sheet5C364DB7AorB 10K
R378 register4rregisterflipflop3andd1sheet5C364DB7B register4rregisterflipflop3andd1sheet5C364DB7AorB 10K
Q150 register4rregisterflipflop3andd1Q register4rregisterflipflop3andd1sheet5C364DB7AorB 0 NPN
R381 adder4Vcc register4rregisterflipflop3andd1sheet5C364DB7A 1K
R380 register4rD3 register4rregisterflipflop3andd1Sheet5C3654CCQr 10K
Q151 register4rregisterflipflop3andd1sheet5C364DB7A register4rregisterflipflop3andd1Sheet5C3654CCQr 0 NPN
R383 adder4Vcc register4rregisterflipflop3andd1sheet5C364DB7B 1K
R382 register4aCLK register4rregisterflipflop3andd1sheet5C366192Qr 10K
Q152 register4rregisterflipflop3andd1sheet5C364DB7B register4rregisterflipflop3andd1sheet5C366192Qr 0 NPN
R385 adder4Vcc register4rregisterflipflop3andd2B 1K
R384 register4rD3 register4rregisterflipflop3notd1Qr 10K
Q153 register4rregisterflipflop3andd2B register4rregisterflipflop3notd1Qr 0 NPN
R387 adder4Vcc register4rregisterflipflop3notd3NQ 1K
R386 register4rregisterflipflop3andd2Q register4rregisterflipflop3notd3Qr 10K
Q154 register4rregisterflipflop3notd3NQ register4rregisterflipflop3notd3Qr 0 NPN
R390 adder4Vcc register4rregisterflipflop3andd2Q 1K
R388 register4rregisterflipflop3andd2sheet5C364DB7A register4rregisterflipflop3andd2sheet5C364DB7AorB 10K
R389 register4rregisterflipflop3andd2sheet5C364DB7B register4rregisterflipflop3andd2sheet5C364DB7AorB 10K
Q155 register4rregisterflipflop3andd2Q register4rregisterflipflop3andd2sheet5C364DB7AorB 0 NPN
R392 adder4Vcc register4rregisterflipflop3andd2sheet5C364DB7A 1K
R391 register4aCLK register4rregisterflipflop3andd2Sheet5C3654CCQr 10K
Q156 register4rregisterflipflop3andd2sheet5C364DB7A register4rregisterflipflop3andd2Sheet5C3654CCQr 0 NPN
R394 adder4Vcc register4rregisterflipflop3andd2sheet5C364DB7B 1K
R393 register4rregisterflipflop3andd2B register4rregisterflipflop3andd2sheet5C366192Qr 10K
Q157 register4rregisterflipflop3andd2sheet5C364DB7B register4rregisterflipflop3andd2sheet5C366192Qr 0 NPN
R397 adder4Vcc register4rQ4 1K
R395 register4rregisterflipflop4notd3NQ register4rregisterflipflop4srlatchdsheet5C3630E6AorB 10K
R396 register4rregisterflipflop4NQ register4rregisterflipflop4srlatchdsheet5C3630E6AorB 10K
Q158 register4rQ4 register4rregisterflipflop4srlatchdsheet5C3630E6AorB 0 NPN
R400 adder4Vcc register4rregisterflipflop4NQ 1K
R398 register4rQ4 register4rregisterflipflop4srlatchdsheet5C3630F6AorB 10K
R399 register4rregisterflipflop4notd2NQ register4rregisterflipflop4srlatchdsheet5C3630F6AorB 10K
Q159 register4rregisterflipflop4NQ register4rregisterflipflop4srlatchdsheet5C3630F6AorB 0 NPN
R402 adder4Vcc register4rregisterflipflop4notd2NQ 1K
R401 register4rregisterflipflop4andd1Q register4rregisterflipflop4notd2Qr 10K
Q160 register4rregisterflipflop4notd2NQ register4rregisterflipflop4notd2Qr 0 NPN
R405 adder4Vcc register4rregisterflipflop4andd1Q 1K
R403 register4rregisterflipflop4andd1sheet5C364DB7A register4rregisterflipflop4andd1sheet5C364DB7AorB 10K
R404 register4rregisterflipflop4andd1sheet5C364DB7B register4rregisterflipflop4andd1sheet5C364DB7AorB 10K
Q161 register4rregisterflipflop4andd1Q register4rregisterflipflop4andd1sheet5C364DB7AorB 0 NPN
R407 adder4Vcc register4rregisterflipflop4andd1sheet5C364DB7A 1K
R406 register4rD4 register4rregisterflipflop4andd1Sheet5C3654CCQr 10K
Q162 register4rregisterflipflop4andd1sheet5C364DB7A register4rregisterflipflop4andd1Sheet5C3654CCQr 0 NPN
R409 adder4Vcc register4rregisterflipflop4andd1sheet5C364DB7B 1K
R408 register4aCLK register4rregisterflipflop4andd1sheet5C366192Qr 10K
Q163 register4rregisterflipflop4andd1sheet5C364DB7B register4rregisterflipflop4andd1sheet5C366192Qr 0 NPN
R411 adder4Vcc register4rregisterflipflop4andd2B 1K
R410 register4rD4 register4rregisterflipflop4notd1Qr 10K
Q164 register4rregisterflipflop4andd2B register4rregisterflipflop4notd1Qr 0 NPN
R413 adder4Vcc register4rregisterflipflop4notd3NQ 1K
R412 register4rregisterflipflop4andd2Q register4rregisterflipflop4notd3Qr 10K
Q165 register4rregisterflipflop4notd3NQ register4rregisterflipflop4notd3Qr 0 NPN
R416 adder4Vcc register4rregisterflipflop4andd2Q 1K
R414 register4rregisterflipflop4andd2sheet5C364DB7A register4rregisterflipflop4andd2sheet5C364DB7AorB 10K
R415 register4rregisterflipflop4andd2sheet5C364DB7B register4rregisterflipflop4andd2sheet5C364DB7AorB 10K
Q166 register4rregisterflipflop4andd2Q register4rregisterflipflop4andd2sheet5C364DB7AorB 0 NPN
R418 adder4Vcc register4rregisterflipflop4andd2sheet5C364DB7A 1K
R417 register4aCLK register4rregisterflipflop4andd2Sheet5C3654CCQr 10K
Q167 register4rregisterflipflop4andd2sheet5C364DB7A register4rregisterflipflop4andd2Sheet5C3654CCQr 0 NPN
R420 adder4Vcc register4rregisterflipflop4andd2sheet5C364DB7B 1K
R419 register4rregisterflipflop4andd2B register4rregisterflipflop4andd2sheet5C366192Qr 10K
Q168 register4rregisterflipflop4andd2sheet5C364DB7B register4rregisterflipflop4andd2sheet5C366192Qr 0 NPN
.op
.dc v1 5 5 1
.print dc i(v1)
.end
