.title KiCad schematic
.op
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V3 and42Vcc 0 dc 5
V1 A1 0 dc 0
V2 A2 0 dc 5
V4 A3 0 dc 0
V5 A4 0 dc 5
V6 B1 0 dc 5
V7 and42B2 0 dc 5
V8 B3 0 dc 5
V9 B4 0 dc 5
R3 and42Vcc and42Q1 1K
R1 and42gateand42and1sheet5C364DB7A and42gateand42and1sheet5C364DB7AorB 10K
R2 and42gateand42and1sheet5C364DB7B and42gateand42and1sheet5C364DB7AorB 10K
Q1 and42Q1 and42gateand42and1sheet5C364DB7AorB 0 NPN
R5 and42Vcc and42gateand42and1sheet5C364DB7A 1K
R4 A1 and42gateand42and1Sheet5C3654CCQr 10K
Q2 and42gateand42and1sheet5C364DB7A and42gateand42and1Sheet5C3654CCQr 0 NPN
R7 and42Vcc and42gateand42and1sheet5C364DB7B 1K
R6 B1 and42gateand42and1sheet5C366192Qr 10K
Q3 and42gateand42and1sheet5C364DB7B and42gateand42and1sheet5C366192Qr 0 NPN
R10 and42Vcc and42Q2 1K
R8 and42gateand42and2sheet5C364DB7A and42gateand42and2sheet5C364DB7AorB 10K
R9 and42gateand42and2sheet5C364DB7B and42gateand42and2sheet5C364DB7AorB 10K
Q4 and42Q2 and42gateand42and2sheet5C364DB7AorB 0 NPN
R12 and42Vcc and42gateand42and2sheet5C364DB7A 1K
R11 A2 and42gateand42and2Sheet5C3654CCQr 10K
Q5 and42gateand42and2sheet5C364DB7A and42gateand42and2Sheet5C3654CCQr 0 NPN
R14 and42Vcc and42gateand42and2sheet5C364DB7B 1K
R13 and42B2 and42gateand42and2sheet5C366192Qr 10K
Q6 and42gateand42and2sheet5C364DB7B and42gateand42and2sheet5C366192Qr 0 NPN
R17 and42Vcc and42Q3 1K
R15 and42gateand42and3sheet5C364DB7A and42gateand42and3sheet5C364DB7AorB 10K
R16 and42gateand42and3sheet5C364DB7B and42gateand42and3sheet5C364DB7AorB 10K
Q7 and42Q3 and42gateand42and3sheet5C364DB7AorB 0 NPN
R19 and42Vcc and42gateand42and3sheet5C364DB7A 1K
R18 A3 and42gateand42and3Sheet5C3654CCQr 10K
Q8 and42gateand42and3sheet5C364DB7A and42gateand42and3Sheet5C3654CCQr 0 NPN
R21 and42Vcc and42gateand42and3sheet5C364DB7B 1K
R20 B3 and42gateand42and3sheet5C366192Qr 10K
Q9 and42gateand42and3sheet5C364DB7B and42gateand42and3sheet5C366192Qr 0 NPN
R24 and42Vcc and42Q4 1K
R22 and42gateand42and4sheet5C364DB7A and42gateand42and4sheet5C364DB7AorB 10K
R23 and42gateand42and4sheet5C364DB7B and42gateand42and4sheet5C364DB7AorB 10K
Q10 and42Q4 and42gateand42and4sheet5C364DB7AorB 0 NPN
R26 and42Vcc and42gateand42and4sheet5C364DB7A 1K
R25 A4 and42gateand42and4Sheet5C3654CCQr 10K
Q11 and42gateand42and4sheet5C364DB7A and42gateand42and4Sheet5C3654CCQr 0 NPN
R28 and42Vcc and42gateand42and4sheet5C364DB7B 1K
R27 B4 and42gateand42and4sheet5C366192Qr 10K
Q12 and42gateand42and4sheet5C364DB7B and42gateand42and4sheet5C366192Qr 0 NPN
.end
