.title KiCad schematic
.op
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V4 adder4Vcc 0 dc 5
V1 A1in 0 dc 5
V2 A2in 0 dc 5
V3 A3in 0 dc 0
V5 A4in 0 dc 0
V6 B1in 0 dc 0
V7 B2in 0 dc 5
V8 B3in 0 dc 0
V9 B4in 0 dc 0
V10 Cinin 0 dc 0
R3 adder4Vcc adder4adder41sheet5C34B00DA 1K
R1 A1in adder4adder41sheet5C34AF27AorB 10K
R2 B1in adder4adder41sheet5C34AF27AorB 10K
Q1 adder4adder41sheet5C34B00DA adder4adder41sheet5C34AF27AorB 0 NPN
R6 adder4Vcc adder4adder41sheet5C34B027A 1K
R4 A1in adder4adder41sheet5C34AFF9AorB 10K
R5 adder4adder41sheet5C34B00DA adder4adder41sheet5C34AFF9AorB 10K
Q2 adder4adder41sheet5C34B027A adder4adder41sheet5C34AFF9AorB 0 NPN
R9 adder4Vcc adder4adder41sheet5C34B027B 1K
R7 adder4adder41sheet5C34B00DA adder4adder41sheet5C34B00DAorB 10K
R8 B1in adder4adder41sheet5C34B00DAorB 10K
Q3 adder4adder41sheet5C34B027B adder4adder41sheet5C34B00DAorB 0 NPN
R12 adder4Vcc adder4adder41sheet5C34B047A 1K
R10 adder4adder41sheet5C34B027A adder4adder41sheet5C34B027AorB 10K
R11 adder4adder41sheet5C34B027B adder4adder41sheet5C34B027AorB 10K
Q4 adder4adder41sheet5C34B047A adder4adder41sheet5C34B027AorB 0 NPN
R15 adder4Vcc adder4adder41sheet5C34B049A 1K
R13 adder4adder41sheet5C34B047A adder4adder41sheet5C34B047AorB 10K
R14 Cinin adder4adder41sheet5C34B047AorB 10K
Q5 adder4adder41sheet5C34B049A adder4adder41sheet5C34B047AorB 0 NPN
R18 adder4Vcc adder4adder41sheet5C34B04AA 1K
R16 adder4adder41sheet5C34B047A adder4adder41sheet5C34B048AorB 10K
R17 adder4adder41sheet5C34B049A adder4adder41sheet5C34B048AorB 10K
Q6 adder4adder41sheet5C34B04AA adder4adder41sheet5C34B048AorB 0 NPN
R21 adder4Vcc adder4adder41sheet5C34B04AB 1K
R19 adder4adder41sheet5C34B049A adder4adder41sheet5C34B049AorB 10K
R20 Cinin adder4adder41sheet5C34B049AorB 10K
Q7 adder4adder41sheet5C34B04AB adder4adder41sheet5C34B049AorB 0 NPN
R24 adder4Vcc adder4S1 1K
R22 adder4adder41sheet5C34B04AA adder4adder41sheet5C34B04AAorB 10K
R23 adder4adder41sheet5C34B04AB adder4adder41sheet5C34B04AAorB 10K
Q8 adder4S1 adder4adder41sheet5C34B04AAorB 0 NPN
R27 adder4Vcc adder4adder42Cin 1K
R25 adder4adder41sheet5C34B049A adder4adder41sheet5C34B0CDAorB 10K
R26 adder4adder41sheet5C34B00DA adder4adder41sheet5C34B0CDAorB 10K
Q9 adder4adder42Cin adder4adder41sheet5C34B0CDAorB 0 NPN
R30 adder4Vcc adder4adder42sheet5C34B00DA 1K
R28 A2in adder4adder42sheet5C34AF27AorB 10K
R29 B2in adder4adder42sheet5C34AF27AorB 10K
Q10 adder4adder42sheet5C34B00DA adder4adder42sheet5C34AF27AorB 0 NPN
R33 adder4Vcc adder4adder42sheet5C34B027A 1K
R31 A2in adder4adder42sheet5C34AFF9AorB 10K
R32 adder4adder42sheet5C34B00DA adder4adder42sheet5C34AFF9AorB 10K
Q11 adder4adder42sheet5C34B027A adder4adder42sheet5C34AFF9AorB 0 NPN
R36 adder4Vcc adder4adder42sheet5C34B027B 1K
R34 adder4adder42sheet5C34B00DA adder4adder42sheet5C34B00DAorB 10K
R35 B2in adder4adder42sheet5C34B00DAorB 10K
Q12 adder4adder42sheet5C34B027B adder4adder42sheet5C34B00DAorB 0 NPN
R39 adder4Vcc adder4adder42sheet5C34B047A 1K
R37 adder4adder42sheet5C34B027A adder4adder42sheet5C34B027AorB 10K
R38 adder4adder42sheet5C34B027B adder4adder42sheet5C34B027AorB 10K
Q13 adder4adder42sheet5C34B047A adder4adder42sheet5C34B027AorB 0 NPN
R42 adder4Vcc adder4adder42sheet5C34B049A 1K
R40 adder4adder42sheet5C34B047A adder4adder42sheet5C34B047AorB 10K
R41 adder4adder42Cin adder4adder42sheet5C34B047AorB 10K
Q14 adder4adder42sheet5C34B049A adder4adder42sheet5C34B047AorB 0 NPN
R45 adder4Vcc adder4adder42sheet5C34B04AA 1K
R43 adder4adder42sheet5C34B047A adder4adder42sheet5C34B048AorB 10K
R44 adder4adder42sheet5C34B049A adder4adder42sheet5C34B048AorB 10K
Q15 adder4adder42sheet5C34B04AA adder4adder42sheet5C34B048AorB 0 NPN
R48 adder4Vcc adder4adder42sheet5C34B04AB 1K
R46 adder4adder42sheet5C34B049A adder4adder42sheet5C34B049AorB 10K
R47 adder4adder42Cin adder4adder42sheet5C34B049AorB 10K
Q16 adder4adder42sheet5C34B04AB adder4adder42sheet5C34B049AorB 0 NPN
R51 adder4Vcc adder4S2 1K
R49 adder4adder42sheet5C34B04AA adder4adder42sheet5C34B04AAorB 10K
R50 adder4adder42sheet5C34B04AB adder4adder42sheet5C34B04AAorB 10K
Q17 adder4S2 adder4adder42sheet5C34B04AAorB 0 NPN
R54 adder4Vcc adder4adder43Cin 1K
R52 adder4adder42sheet5C34B049A adder4adder42sheet5C34B0CDAorB 10K
R53 adder4adder42sheet5C34B00DA adder4adder42sheet5C34B0CDAorB 10K
Q18 adder4adder43Cin adder4adder42sheet5C34B0CDAorB 0 NPN
R57 adder4Vcc adder4adder43sheet5C34B00DA 1K
R55 A3in adder4adder43sheet5C34AF27AorB 10K
R56 B3in adder4adder43sheet5C34AF27AorB 10K
Q19 adder4adder43sheet5C34B00DA adder4adder43sheet5C34AF27AorB 0 NPN
R60 adder4Vcc adder4adder43sheet5C34B027A 1K
R58 A3in adder4adder43sheet5C34AFF9AorB 10K
R59 adder4adder43sheet5C34B00DA adder4adder43sheet5C34AFF9AorB 10K
Q20 adder4adder43sheet5C34B027A adder4adder43sheet5C34AFF9AorB 0 NPN
R63 adder4Vcc adder4adder43sheet5C34B027B 1K
R61 adder4adder43sheet5C34B00DA adder4adder43sheet5C34B00DAorB 10K
R62 B3in adder4adder43sheet5C34B00DAorB 10K
Q21 adder4adder43sheet5C34B027B adder4adder43sheet5C34B00DAorB 0 NPN
R66 adder4Vcc adder4adder43sheet5C34B047A 1K
R64 adder4adder43sheet5C34B027A adder4adder43sheet5C34B027AorB 10K
R65 adder4adder43sheet5C34B027B adder4adder43sheet5C34B027AorB 10K
Q22 adder4adder43sheet5C34B047A adder4adder43sheet5C34B027AorB 0 NPN
R69 adder4Vcc adder4adder43sheet5C34B049A 1K
R67 adder4adder43sheet5C34B047A adder4adder43sheet5C34B047AorB 10K
R68 adder4adder43Cin adder4adder43sheet5C34B047AorB 10K
Q23 adder4adder43sheet5C34B049A adder4adder43sheet5C34B047AorB 0 NPN
R72 adder4Vcc adder4adder43sheet5C34B04AA 1K
R70 adder4adder43sheet5C34B047A adder4adder43sheet5C34B048AorB 10K
R71 adder4adder43sheet5C34B049A adder4adder43sheet5C34B048AorB 10K
Q24 adder4adder43sheet5C34B04AA adder4adder43sheet5C34B048AorB 0 NPN
R75 adder4Vcc adder4adder43sheet5C34B04AB 1K
R73 adder4adder43sheet5C34B049A adder4adder43sheet5C34B049AorB 10K
R74 adder4adder43Cin adder4adder43sheet5C34B049AorB 10K
Q25 adder4adder43sheet5C34B04AB adder4adder43sheet5C34B049AorB 0 NPN
R78 adder4Vcc adder4S3 1K
R76 adder4adder43sheet5C34B04AA adder4adder43sheet5C34B04AAorB 10K
R77 adder4adder43sheet5C34B04AB adder4adder43sheet5C34B04AAorB 10K
Q26 adder4S3 adder4adder43sheet5C34B04AAorB 0 NPN
R81 adder4Vcc adder4adder44Cin 1K
R79 adder4adder43sheet5C34B049A adder4adder43sheet5C34B0CDAorB 10K
R80 adder4adder43sheet5C34B00DA adder4adder43sheet5C34B0CDAorB 10K
Q27 adder4adder44Cin adder4adder43sheet5C34B0CDAorB 0 NPN
R84 adder4Vcc adder4adder44sheet5C34B00DA 1K
R82 A4in adder4adder44sheet5C34AF27AorB 10K
R83 B4in adder4adder44sheet5C34AF27AorB 10K
Q28 adder4adder44sheet5C34B00DA adder4adder44sheet5C34AF27AorB 0 NPN
R87 adder4Vcc adder4adder44sheet5C34B027A 1K
R85 A4in adder4adder44sheet5C34AFF9AorB 10K
R86 adder4adder44sheet5C34B00DA adder4adder44sheet5C34AFF9AorB 10K
Q29 adder4adder44sheet5C34B027A adder4adder44sheet5C34AFF9AorB 0 NPN
R90 adder4Vcc adder4adder44sheet5C34B027B 1K
R88 adder4adder44sheet5C34B00DA adder4adder44sheet5C34B00DAorB 10K
R89 B4in adder4adder44sheet5C34B00DAorB 10K
Q30 adder4adder44sheet5C34B027B adder4adder44sheet5C34B00DAorB 0 NPN
R93 adder4Vcc adder4adder44sheet5C34B047A 1K
R91 adder4adder44sheet5C34B027A adder4adder44sheet5C34B027AorB 10K
R92 adder4adder44sheet5C34B027B adder4adder44sheet5C34B027AorB 10K
Q31 adder4adder44sheet5C34B047A adder4adder44sheet5C34B027AorB 0 NPN
R96 adder4Vcc adder4adder44sheet5C34B049A 1K
R94 adder4adder44sheet5C34B047A adder4adder44sheet5C34B047AorB 10K
R95 adder4adder44Cin adder4adder44sheet5C34B047AorB 10K
Q32 adder4adder44sheet5C34B049A adder4adder44sheet5C34B047AorB 0 NPN
R99 adder4Vcc adder4adder44sheet5C34B04AA 1K
R97 adder4adder44sheet5C34B047A adder4adder44sheet5C34B048AorB 10K
R98 adder4adder44sheet5C34B049A adder4adder44sheet5C34B048AorB 10K
Q33 adder4adder44sheet5C34B04AA adder4adder44sheet5C34B048AorB 0 NPN
R102 adder4Vcc adder4adder44sheet5C34B04AB 1K
R100 adder4adder44sheet5C34B049A adder4adder44sheet5C34B049AorB 10K
R101 adder4adder44Cin adder4adder44sheet5C34B049AorB 10K
Q34 adder4adder44sheet5C34B04AB adder4adder44sheet5C34B049AorB 0 NPN
R105 adder4Vcc adder4S4 1K
R103 adder4adder44sheet5C34B04AA adder4adder44sheet5C34B04AAorB 10K
R104 adder4adder44sheet5C34B04AB adder4adder44sheet5C34B04AAorB 10K
Q35 adder4S4 adder4adder44sheet5C34B04AAorB 0 NPN
R108 adder4Vcc adder4Cout 1K
R106 adder4adder44sheet5C34B049A adder4adder44sheet5C34B0CDAorB 10K
R107 adder4adder44sheet5C34B00DA adder4adder44sheet5C34B0CDAorB 10K
Q36 adder4Cout adder4adder44sheet5C34B0CDAorB 0 NPN
.end
