.title KiCad schematic
V1 /not/Vcc 0 dc 5
V2 /Qin 0 dc 5
R2 /not/Vcc /Q 1K
R1 /Qin /not/Qr 10K
Q1 /Q /not/Qr 0 NPN
.end
