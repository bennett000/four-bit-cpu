.title KiCad schematic
* .op
.tran 1ns 500ns
.print tran v(aluz1) v(aluz2) v(aluz3) v(aluz4)
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V14 aluVcc 0 dc 5
V1 B1in 0 dc 0
V2 B2in 0 dc 5
V3 B3in 0 dc 0
V5 B4in 0 dc 0
V10 A1in 0 dc 5
V11 A2in 0 dc 5
V12 A3in 0 dc 0
V13 A4in 0 dc 0
V4 S1 0 dc 0
V6 S2 0 dc 0
V7 S3 0 dc 0
V8 S4 0 dc 0
V9 S0 0 dc 0
R2 aluVcc alualureplicate141replicate14buffer1buffernot1NQ 1K
R1 alualureplicate141A alualureplicate141replicate14buffer1buffernot1Qr 10K
Q1 alualureplicate141replicate14buffer1buffernot1NQ alualureplicate141replicate14buffer1buffernot1Qr 0 NPN
R4 aluVcc alualuand41A1 1K
R3 alualureplicate141replicate14buffer1buffernot1NQ alualureplicate141replicate14buffer1buffernot2Qr 10K
Q2 alualuand41A1 alualureplicate141replicate14buffer1buffernot2Qr 0 NPN
R6 aluVcc alualureplicate141replicate14buffer2buffernot1NQ 1K
R5 alualureplicate141A alualureplicate141replicate14buffer2buffernot1Qr 10K
Q3 alualureplicate141replicate14buffer2buffernot1NQ alualureplicate141replicate14buffer2buffernot1Qr 0 NPN
R8 aluVcc alualuand41A2 1K
R7 alualureplicate141replicate14buffer2buffernot1NQ alualureplicate141replicate14buffer2buffernot2Qr 10K
Q4 alualuand41A2 alualureplicate141replicate14buffer2buffernot2Qr 0 NPN
R10 aluVcc alualureplicate141replicate14buffer3buffernot1NQ 1K
R9 alualureplicate141A alualureplicate141replicate14buffer3buffernot1Qr 10K
Q5 alualureplicate141replicate14buffer3buffernot1NQ alualureplicate141replicate14buffer3buffernot1Qr 0 NPN
R12 aluVcc alualuand41A3 1K
R11 alualureplicate141replicate14buffer3buffernot1NQ alualureplicate141replicate14buffer3buffernot2Qr 10K
Q6 alualuand41A3 alualureplicate141replicate14buffer3buffernot2Qr 0 NPN
R14 aluVcc alualureplicate141replicate14buffer4buffernot1NQ 1K
R13 alualureplicate141A alualureplicate141replicate14buffer4buffernot1Qr 10K
Q7 alualureplicate141replicate14buffer4buffernot1NQ alualureplicate141replicate14buffer4buffernot1Qr 0 NPN
R16 aluVcc alualuand41A4 1K
R15 alualureplicate141replicate14buffer4buffernot1NQ alualureplicate141replicate14buffer4buffernot2Qr 10K
Q8 alualuand41A4 alualureplicate141replicate14buffer4buffernot2Qr 0 NPN
R19 aluVcc alualumux4411B1 1K
R17 alualuand42gateand42and1sheet5C364DB7A alualuand42gateand42and1sheet5C364DB7AorB 10K
R18 alualuand42gateand42and1sheet5C364DB7B alualuand42gateand42and1sheet5C364DB7AorB 10K
Q9 alualumux4411B1 alualuand42gateand42and1sheet5C364DB7AorB 0 NPN
R21 aluVcc alualuand42gateand42and1sheet5C364DB7A 1K
R20 A1in alualuand42gateand42and1Sheet5C3654CCQr 10K
Q10 alualuand42gateand42and1sheet5C364DB7A alualuand42gateand42and1Sheet5C3654CCQr 0 NPN
R23 aluVcc alualuand42gateand42and1sheet5C364DB7B 1K
R22 B1in alualuand42gateand42and1sheet5C366192Qr 10K
Q11 alualuand42gateand42and1sheet5C364DB7B alualuand42gateand42and1sheet5C366192Qr 0 NPN
R26 aluVcc alualumux4411B2 1K
R24 alualuand42gateand42and2sheet5C364DB7A alualuand42gateand42and2sheet5C364DB7AorB 10K
R25 alualuand42gateand42and2sheet5C364DB7B alualuand42gateand42and2sheet5C364DB7AorB 10K
Q12 alualumux4411B2 alualuand42gateand42and2sheet5C364DB7AorB 0 NPN
R28 aluVcc alualuand42gateand42and2sheet5C364DB7A 1K
R27 A2in alualuand42gateand42and2Sheet5C3654CCQr 10K
Q13 alualuand42gateand42and2sheet5C364DB7A alualuand42gateand42and2Sheet5C3654CCQr 0 NPN
R30 aluVcc alualuand42gateand42and2sheet5C364DB7B 1K
R29 B2in alualuand42gateand42and2sheet5C366192Qr 10K
Q14 alualuand42gateand42and2sheet5C364DB7B alualuand42gateand42and2sheet5C366192Qr 0 NPN
R33 aluVcc alualumux4411B3 1K
R31 alualuand42gateand42and3sheet5C364DB7A alualuand42gateand42and3sheet5C364DB7AorB 10K
R32 alualuand42gateand42and3sheet5C364DB7B alualuand42gateand42and3sheet5C364DB7AorB 10K
Q15 alualumux4411B3 alualuand42gateand42and3sheet5C364DB7AorB 0 NPN
R35 aluVcc alualuand42gateand42and3sheet5C364DB7A 1K
R34 A3in alualuand42gateand42and3Sheet5C3654CCQr 10K
Q16 alualuand42gateand42and3sheet5C364DB7A alualuand42gateand42and3Sheet5C3654CCQr 0 NPN
R37 aluVcc alualuand42gateand42and3sheet5C364DB7B 1K
R36 B3in alualuand42gateand42and3sheet5C366192Qr 10K
Q17 alualuand42gateand42and3sheet5C364DB7B alualuand42gateand42and3sheet5C366192Qr 0 NPN
R40 aluVcc alualumux4411B4 1K
R38 alualuand42gateand42and4sheet5C364DB7A alualuand42gateand42and4sheet5C364DB7AorB 10K
R39 alualuand42gateand42and4sheet5C364DB7B alualuand42gateand42and4sheet5C364DB7AorB 10K
Q18 alualumux4411B4 alualuand42gateand42and4sheet5C364DB7AorB 0 NPN
R42 aluVcc alualuand42gateand42and4sheet5C364DB7A 1K
R41 A4in alualuand42gateand42and4Sheet5C3654CCQr 10K
Q19 alualuand42gateand42and4sheet5C364DB7A alualuand42gateand42and4Sheet5C3654CCQr 0 NPN
R44 aluVcc alualuand42gateand42and4sheet5C364DB7B 1K
R43 B4in alualuand42gateand42and4sheet5C366192Qr 10K
Q20 alualuand42gateand42and4sheet5C364DB7B alualuand42gateand42and4sheet5C366192Qr 0 NPN
R47 aluVcc alualubitwiseinv1bitwiseinvxor21xor2nor2B 1K
R45 S4 alualubitwiseinv1bitwiseinvxor21xor2nor1AorB 10K
R46 B1in alualubitwiseinv1bitwiseinvxor21xor2nor1AorB 10K
Q21 alualubitwiseinv1bitwiseinvxor21xor2nor2B alualubitwiseinv1bitwiseinvxor21xor2nor1AorB 0 NPN
R50 aluVcc alualubitwiseinv1bitwiseinvxor21xor2nor2A 1K
R48 alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7AorB 10K
R49 alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7AorB 10K
Q22 alualubitwiseinv1bitwiseinvxor21xor2nor2A alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7AorB 0 NPN
R52 aluVcc alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7A 1K
R51 S4 alualubitwiseinv1bitwiseinvxor21xor2and1Sheet5C3654CCQr 10K
Q23 alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor21xor2and1Sheet5C3654CCQr 0 NPN
R54 aluVcc alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7B 1K
R53 B1in alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C366192Qr 10K
Q24 alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor21xor2and1sheet5C366192Qr 0 NPN
R57 aluVcc alualuand41B1 1K
R55 alualubitwiseinv1bitwiseinvxor21xor2nor2A alualubitwiseinv1bitwiseinvxor21xor2nor2AorB 10K
R56 alualubitwiseinv1bitwiseinvxor21xor2nor2B alualubitwiseinv1bitwiseinvxor21xor2nor2AorB 10K
Q25 alualuand41B1 alualubitwiseinv1bitwiseinvxor21xor2nor2AorB 0 NPN
R60 aluVcc alualubitwiseinv1bitwiseinvxor22xor2nor2B 1K
R58 S4 alualubitwiseinv1bitwiseinvxor22xor2nor1AorB 10K
R59 B2in alualubitwiseinv1bitwiseinvxor22xor2nor1AorB 10K
Q26 alualubitwiseinv1bitwiseinvxor22xor2nor2B alualubitwiseinv1bitwiseinvxor22xor2nor1AorB 0 NPN
R63 aluVcc alualubitwiseinv1bitwiseinvxor22xor2nor2A 1K
R61 alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7AorB 10K
R62 alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7AorB 10K
Q27 alualubitwiseinv1bitwiseinvxor22xor2nor2A alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7AorB 0 NPN
R65 aluVcc alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7A 1K
R64 S4 alualubitwiseinv1bitwiseinvxor22xor2and1Sheet5C3654CCQr 10K
Q28 alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor22xor2and1Sheet5C3654CCQr 0 NPN
R67 aluVcc alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7B 1K
R66 B2in alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C366192Qr 10K
Q29 alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor22xor2and1sheet5C366192Qr 0 NPN
R70 aluVcc alualuand41B2 1K
R68 alualubitwiseinv1bitwiseinvxor22xor2nor2A alualubitwiseinv1bitwiseinvxor22xor2nor2AorB 10K
R69 alualubitwiseinv1bitwiseinvxor22xor2nor2B alualubitwiseinv1bitwiseinvxor22xor2nor2AorB 10K
Q30 alualuand41B2 alualubitwiseinv1bitwiseinvxor22xor2nor2AorB 0 NPN
R73 aluVcc alualubitwiseinv1bitwiseinvxor23xor2nor2B 1K
R71 S4 alualubitwiseinv1bitwiseinvxor23xor2nor1AorB 10K
R72 B3in alualubitwiseinv1bitwiseinvxor23xor2nor1AorB 10K
Q31 alualubitwiseinv1bitwiseinvxor23xor2nor2B alualubitwiseinv1bitwiseinvxor23xor2nor1AorB 0 NPN
R76 aluVcc alualubitwiseinv1bitwiseinvxor23xor2nor2A 1K
R74 alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7AorB 10K
R75 alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7AorB 10K
Q32 alualubitwiseinv1bitwiseinvxor23xor2nor2A alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7AorB 0 NPN
R78 aluVcc alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7A 1K
R77 S4 alualubitwiseinv1bitwiseinvxor23xor2and1Sheet5C3654CCQr 10K
Q33 alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor23xor2and1Sheet5C3654CCQr 0 NPN
R80 aluVcc alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7B 1K
R79 B3in alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C366192Qr 10K
Q34 alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor23xor2and1sheet5C366192Qr 0 NPN
R83 aluVcc alualuand41B3 1K
R81 alualubitwiseinv1bitwiseinvxor23xor2nor2A alualubitwiseinv1bitwiseinvxor23xor2nor2AorB 10K
R82 alualubitwiseinv1bitwiseinvxor23xor2nor2B alualubitwiseinv1bitwiseinvxor23xor2nor2AorB 10K
Q35 alualuand41B3 alualubitwiseinv1bitwiseinvxor23xor2nor2AorB 0 NPN
R86 aluVcc alualubitwiseinv1bitwiseinvxor24xor2nor2B 1K
R84 S4 alualubitwiseinv1bitwiseinvxor24xor2nor1AorB 10K
R85 B4in alualubitwiseinv1bitwiseinvxor24xor2nor1AorB 10K
Q36 alualubitwiseinv1bitwiseinvxor24xor2nor2B alualubitwiseinv1bitwiseinvxor24xor2nor1AorB 0 NPN
R89 aluVcc alualubitwiseinv1bitwiseinvxor24xor2nor2A 1K
R87 alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7AorB 10K
R88 alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7AorB 10K
Q37 alualubitwiseinv1bitwiseinvxor24xor2nor2A alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7AorB 0 NPN
R91 aluVcc alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7A 1K
R90 S4 alualubitwiseinv1bitwiseinvxor24xor2and1Sheet5C3654CCQr 10K
Q38 alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7A alualubitwiseinv1bitwiseinvxor24xor2and1Sheet5C3654CCQr 0 NPN
R93 aluVcc alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7B 1K
R92 B4in alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C366192Qr 10K
Q39 alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C364DB7B alualubitwiseinv1bitwiseinvxor24xor2and1sheet5C366192Qr 0 NPN
R96 aluVcc alualuand41B4 1K
R94 alualubitwiseinv1bitwiseinvxor24xor2nor2A alualubitwiseinv1bitwiseinvxor24xor2nor2AorB 10K
R95 alualubitwiseinv1bitwiseinvxor24xor2nor2B alualubitwiseinv1bitwiseinvxor24xor2nor2AorB 10K
Q40 alualuand41B4 alualubitwiseinv1bitwiseinvxor24xor2nor2AorB 0 NPN
R98 aluVcc alualumux4411multiplexer441mux4213A1 1K
R97 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornot1Qr 10K
Q41 alualumux4411multiplexer441mux4213A1 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R101 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornor1Q 1K
R99 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornor1AorB 10K
R100 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornor1AorB 10K
Q42 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R104 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1A 1K
R102 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R103 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q43 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R106 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R105 aluAdderS1 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q44 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R108 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R107 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q45 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R111 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1B 1K
R109 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R110 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q46 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R113 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R112 S1 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q47 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R115 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R114 alualumux4411B1 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q48 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R117 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1B 1K
R116 S1 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21not1Qr 10K
Q49 alualumux4411multiplexer441mux4211multiplexer421mux1211mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1211mux21not1Qr 0 NPN
R119 aluVcc alualumux4411multiplexer441mux4213A2 1K
R118 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornot1Qr 10K
Q50 alualumux4411multiplexer441mux4213A2 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R122 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornor1Q 1K
R120 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornor1AorB 10K
R121 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornor1AorB 10K
Q51 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R125 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1A 1K
R123 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R124 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q52 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R127 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R126 aluAdderS1 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q53 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R129 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R128 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q54 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R132 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1B 1K
R130 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R131 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q55 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R134 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R133 S1 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q56 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R136 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R135 alualumux4411B2 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q57 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R138 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1B 1K
R137 S1 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21not1Qr 10K
Q58 alualumux4411multiplexer441mux4211multiplexer421mux1212mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1212mux21not1Qr 0 NPN
R140 aluVcc alualumux4411multiplexer441mux4213A3 1K
R139 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornot1Qr 10K
Q59 alualumux4411multiplexer441mux4213A3 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R143 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornor1Q 1K
R141 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornor1AorB 10K
R142 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornor1AorB 10K
Q60 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R146 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1A 1K
R144 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R145 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q61 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R148 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R147 aluAdderS3 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q62 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R150 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R149 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q63 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R153 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1B 1K
R151 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R152 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q64 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R155 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R154 S1 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q65 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R157 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R156 alualumux4411B3 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q66 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R159 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1B 1K
R158 S1 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21not1Qr 10K
Q67 alualumux4411multiplexer441mux4211multiplexer421mux1213mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1213mux21not1Qr 0 NPN
R161 aluVcc alualumux4411multiplexer441mux4213A4 1K
R160 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornot1Qr 10K
Q68 alualumux4411multiplexer441mux4213A4 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R164 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornor1Q 1K
R162 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornor1AorB 10K
R163 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornor1AorB 10K
Q69 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornor1Q alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R167 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1A 1K
R165 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R166 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q70 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1A alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R169 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R168 aluAdderS4 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q71 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R171 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R170 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q72 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R174 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1B 1K
R172 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R173 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q73 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21or1B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R176 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R175 S1 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q74 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R178 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R177 alualumux4411B4 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q75 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R180 aluVcc alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1B 1K
R179 S1 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21not1Qr 10K
Q76 alualumux4411multiplexer441mux4211multiplexer421mux1214mux21and1B alualumux4411multiplexer441mux4211multiplexer421mux1214mux21not1Qr 0 NPN
R182 aluVcc alualumux4411multiplexer441mux4213B1 1K
R181 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornot1Qr 10K
Q77 alualumux4411multiplexer441mux4213B1 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R185 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornor1Q 1K
R183 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornor1AorB 10K
R184 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornor1AorB 10K
Q78 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R188 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1A 1K
R186 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R187 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q79 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R190 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R189 A1in alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q80 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R192 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R191 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q81 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R195 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1B 1K
R193 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R194 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q82 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R197 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R196 S1 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q83 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R199 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R198 B1in alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q84 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R201 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1B 1K
R200 S1 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21not1Qr 10K
Q85 alualumux4411multiplexer441mux4212multiplexer421mux1211mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1211mux21not1Qr 0 NPN
R203 aluVcc alualumux4411multiplexer441mux4213B2 1K
R202 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornot1Qr 10K
Q86 alualumux4411multiplexer441mux4213B2 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R206 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornor1Q 1K
R204 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornor1AorB 10K
R205 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornor1AorB 10K
Q87 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R209 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1A 1K
R207 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R208 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q88 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R211 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R210 A2in alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q89 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R213 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R212 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q90 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R216 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1B 1K
R214 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R215 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q91 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R218 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R217 S1 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q92 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R220 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R219 B2in alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q93 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R222 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1B 1K
R221 S1 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21not1Qr 10K
Q94 alualumux4411multiplexer441mux4212multiplexer421mux1212mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1212mux21not1Qr 0 NPN
R224 aluVcc alualumux4411multiplexer441mux4213B3 1K
R223 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornot1Qr 10K
Q95 alualumux4411multiplexer441mux4213B3 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R227 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornor1Q 1K
R225 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornor1AorB 10K
R226 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornor1AorB 10K
Q96 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R230 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1A 1K
R228 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R229 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q97 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R232 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R231 A3in alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q98 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R234 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R233 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q99 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R237 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1B 1K
R235 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R236 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q100 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R239 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R238 S1 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q101 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R241 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R240 B3in alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q102 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R243 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1B 1K
R242 S1 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21not1Qr 10K
Q103 alualumux4411multiplexer441mux4212multiplexer421mux1213mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1213mux21not1Qr 0 NPN
R245 aluVcc alualumux4411multiplexer441mux4213B4 1K
R244 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornot1Qr 10K
Q104 alualumux4411multiplexer441mux4213B4 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R248 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornor1Q 1K
R246 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornor1AorB 10K
R247 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornor1AorB 10K
Q105 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornor1Q alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R251 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1A 1K
R249 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R250 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q106 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1A alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R253 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R252 A4in alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q107 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R255 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R254 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q108 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R258 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1B 1K
R256 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R257 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q109 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21or1B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R260 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R259 S1 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q110 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R262 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R261 B4in alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q111 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R264 aluVcc alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1B 1K
R263 S1 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21not1Qr 10K
Q112 alualumux4411multiplexer441mux4212multiplexer421mux1214mux21and1B alualumux4411multiplexer441mux4212multiplexer421mux1214mux21not1Qr 0 NPN
R266 aluVcc aluZ1 1K
R265 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornot1Qr 10K
Q113 aluZ1 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R269 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornor1Q 1K
R267 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornor1AorB 10K
R268 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornor1AorB 10K
Q114 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R272 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1A 1K
R270 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R271 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q115 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R274 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R273 alualumux4411multiplexer441mux4213A1 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q116 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R276 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R275 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q117 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R279 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1B 1K
R277 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R278 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q118 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R281 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R280 S2 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q119 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R283 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R282 alualumux4411multiplexer441mux4213B1 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q120 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R285 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1B 1K
R284 S2 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21not1Qr 10K
Q121 alualumux4411multiplexer441mux4213multiplexer421mux1211mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1211mux21not1Qr 0 NPN
R287 aluVcc aluZ2 1K
R286 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornot1Qr 10K
Q122 aluZ2 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R290 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornor1Q 1K
R288 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornor1AorB 10K
R289 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornor1AorB 10K
Q123 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R293 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1A 1K
R291 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R292 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q124 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R295 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R294 alualumux4411multiplexer441mux4213A2 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q125 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R297 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R296 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q126 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R300 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1B 1K
R298 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R299 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q127 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R302 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R301 S2 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q128 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R304 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R303 alualumux4411multiplexer441mux4213B2 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q129 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R306 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1B 1K
R305 S2 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21not1Qr 10K
Q130 alualumux4411multiplexer441mux4213multiplexer421mux1212mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1212mux21not1Qr 0 NPN
R308 aluVcc aluZ3 1K
R307 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornot1Qr 10K
Q131 aluZ3 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R311 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornor1Q 1K
R309 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornor1AorB 10K
R310 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornor1AorB 10K
Q132 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R314 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1A 1K
R312 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R313 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q133 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R316 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R315 alualumux4411multiplexer441mux4213A3 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q134 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R318 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R317 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q135 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R321 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1B 1K
R319 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R320 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q136 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R323 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R322 S2 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q137 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R325 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R324 alualumux4411multiplexer441mux4213B3 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q138 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R327 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1B 1K
R326 S2 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21not1Qr 10K
Q139 alualumux4411multiplexer441mux4213multiplexer421mux1213mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1213mux21not1Qr 0 NPN
R329 aluVcc aluZ4 1K
R328 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornot1Qr 10K
Q140 aluZ4 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R332 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornor1Q 1K
R330 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornor1AorB 10K
R331 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornor1AorB 10K
Q141 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornor1Q alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R335 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1A 1K
R333 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R334 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q142 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1A alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R337 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R336 alualumux4411multiplexer441mux4213A4 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q143 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R339 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R338 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q144 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R342 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1B 1K
R340 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R341 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q145 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21or1B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R344 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R343 S2 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q146 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7A alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R346 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R345 alualumux4411multiplexer441mux4213B4 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q147 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C364DB7B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R348 aluVcc alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1B 1K
R347 S2 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21not1Qr 10K
Q148 alualumux4411multiplexer441mux4213multiplexer421mux1214mux21and1B alualumux4411multiplexer441mux4213multiplexer421mux1214mux21not1Qr 0 NPN
R351 aluVcc alualuadder41adder41sheet5C34B00DA 1K
R349 A1in alualuadder41adder41sheet5C34AF27AorB 10K
R350 aluAdderB1in alualuadder41adder41sheet5C34AF27AorB 10K
Q149 alualuadder41adder41sheet5C34B00DA alualuadder41adder41sheet5C34AF27AorB 0 NPN
R354 aluVcc alualuadder41adder41sheet5C34B027A 1K
R352 A1in alualuadder41adder41sheet5C34AFF9AorB 10K
R353 alualuadder41adder41sheet5C34B00DA alualuadder41adder41sheet5C34AFF9AorB 10K
Q150 alualuadder41adder41sheet5C34B027A alualuadder41adder41sheet5C34AFF9AorB 0 NPN
R357 aluVcc alualuadder41adder41sheet5C34B027B 1K
R355 alualuadder41adder41sheet5C34B00DA alualuadder41adder41sheet5C34B00DAorB 10K
R356 aluAdderB1in alualuadder41adder41sheet5C34B00DAorB 10K
Q151 alualuadder41adder41sheet5C34B027B alualuadder41adder41sheet5C34B00DAorB 0 NPN
R360 aluVcc alualuadder41adder41sheet5C34B047A 1K
R358 alualuadder41adder41sheet5C34B027A alualuadder41adder41sheet5C34B027AorB 10K
R359 alualuadder41adder41sheet5C34B027B alualuadder41adder41sheet5C34B027AorB 10K
Q152 alualuadder41adder41sheet5C34B047A alualuadder41adder41sheet5C34B027AorB 0 NPN
R363 aluVcc alualuadder41adder41sheet5C34B049A 1K
R361 alualuadder41adder41sheet5C34B047A alualuadder41adder41sheet5C34B047AorB 10K
R362 S3 alualuadder41adder41sheet5C34B047AorB 10K
Q153 alualuadder41adder41sheet5C34B049A alualuadder41adder41sheet5C34B047AorB 0 NPN
R366 aluVcc alualuadder41adder41sheet5C34B04AA 1K
R364 alualuadder41adder41sheet5C34B047A alualuadder41adder41sheet5C34B048AorB 10K
R365 alualuadder41adder41sheet5C34B049A alualuadder41adder41sheet5C34B048AorB 10K
Q154 alualuadder41adder41sheet5C34B04AA alualuadder41adder41sheet5C34B048AorB 0 NPN
R369 aluVcc alualuadder41adder41sheet5C34B04AB 1K
R367 alualuadder41adder41sheet5C34B049A alualuadder41adder41sheet5C34B049AorB 10K
R368 S3 alualuadder41adder41sheet5C34B049AorB 10K
Q155 alualuadder41adder41sheet5C34B04AB alualuadder41adder41sheet5C34B049AorB 0 NPN
R372 aluVcc aluAdderS1 1K
R370 alualuadder41adder41sheet5C34B04AA alualuadder41adder41sheet5C34B04AAorB 10K
R371 alualuadder41adder41sheet5C34B04AB alualuadder41adder41sheet5C34B04AAorB 10K
Q156 aluAdderS1 alualuadder41adder41sheet5C34B04AAorB 0 NPN
R375 aluVcc alualuadder41adder42Cin 1K
R373 alualuadder41adder41sheet5C34B049A alualuadder41adder41sheet5C34B0CDAorB 10K
R374 alualuadder41adder41sheet5C34B00DA alualuadder41adder41sheet5C34B0CDAorB 10K
Q157 alualuadder41adder42Cin alualuadder41adder41sheet5C34B0CDAorB 0 NPN
R378 aluVcc alualuadder41adder42sheet5C34B00DA 1K
R376 A2in alualuadder41adder42sheet5C34AF27AorB 10K
R377 aluAdderB2in alualuadder41adder42sheet5C34AF27AorB 10K
Q158 alualuadder41adder42sheet5C34B00DA alualuadder41adder42sheet5C34AF27AorB 0 NPN
R381 aluVcc alualuadder41adder42sheet5C34B027A 1K
R379 A2in alualuadder41adder42sheet5C34AFF9AorB 10K
R380 alualuadder41adder42sheet5C34B00DA alualuadder41adder42sheet5C34AFF9AorB 10K
Q159 alualuadder41adder42sheet5C34B027A alualuadder41adder42sheet5C34AFF9AorB 0 NPN
R384 aluVcc alualuadder41adder42sheet5C34B027B 1K
R382 alualuadder41adder42sheet5C34B00DA alualuadder41adder42sheet5C34B00DAorB 10K
R383 aluAdderB2in alualuadder41adder42sheet5C34B00DAorB 10K
Q160 alualuadder41adder42sheet5C34B027B alualuadder41adder42sheet5C34B00DAorB 0 NPN
R387 aluVcc alualuadder41adder42sheet5C34B047A 1K
R385 alualuadder41adder42sheet5C34B027A alualuadder41adder42sheet5C34B027AorB 10K
R386 alualuadder41adder42sheet5C34B027B alualuadder41adder42sheet5C34B027AorB 10K
Q161 alualuadder41adder42sheet5C34B047A alualuadder41adder42sheet5C34B027AorB 0 NPN
R390 aluVcc alualuadder41adder42sheet5C34B049A 1K
R388 alualuadder41adder42sheet5C34B047A alualuadder41adder42sheet5C34B047AorB 10K
R389 alualuadder41adder42Cin alualuadder41adder42sheet5C34B047AorB 10K
Q162 alualuadder41adder42sheet5C34B049A alualuadder41adder42sheet5C34B047AorB 0 NPN
R393 aluVcc alualuadder41adder42sheet5C34B04AA 1K
R391 alualuadder41adder42sheet5C34B047A alualuadder41adder42sheet5C34B048AorB 10K
R392 alualuadder41adder42sheet5C34B049A alualuadder41adder42sheet5C34B048AorB 10K
Q163 alualuadder41adder42sheet5C34B04AA alualuadder41adder42sheet5C34B048AorB 0 NPN
R396 aluVcc alualuadder41adder42sheet5C34B04AB 1K
R394 alualuadder41adder42sheet5C34B049A alualuadder41adder42sheet5C34B049AorB 10K
R395 alualuadder41adder42Cin alualuadder41adder42sheet5C34B049AorB 10K
Q164 alualuadder41adder42sheet5C34B04AB alualuadder41adder42sheet5C34B049AorB 0 NPN
R399 aluVcc aluAdderS1 1K
R397 alualuadder41adder42sheet5C34B04AA alualuadder41adder42sheet5C34B04AAorB 10K
R398 alualuadder41adder42sheet5C34B04AB alualuadder41adder42sheet5C34B04AAorB 10K
Q165 aluAdderS1 alualuadder41adder42sheet5C34B04AAorB 0 NPN
R402 aluVcc alualuadder41adder43Cin 1K
R400 alualuadder41adder42sheet5C34B049A alualuadder41adder42sheet5C34B0CDAorB 10K
R401 alualuadder41adder42sheet5C34B00DA alualuadder41adder42sheet5C34B0CDAorB 10K
Q166 alualuadder41adder43Cin alualuadder41adder42sheet5C34B0CDAorB 0 NPN
R405 aluVcc alualuadder41adder43sheet5C34B00DA 1K
R403 A3in alualuadder41adder43sheet5C34AF27AorB 10K
R404 aluAdderB3in alualuadder41adder43sheet5C34AF27AorB 10K
Q167 alualuadder41adder43sheet5C34B00DA alualuadder41adder43sheet5C34AF27AorB 0 NPN
R408 aluVcc alualuadder41adder43sheet5C34B027A 1K
R406 A3in alualuadder41adder43sheet5C34AFF9AorB 10K
R407 alualuadder41adder43sheet5C34B00DA alualuadder41adder43sheet5C34AFF9AorB 10K
Q168 alualuadder41adder43sheet5C34B027A alualuadder41adder43sheet5C34AFF9AorB 0 NPN
R411 aluVcc alualuadder41adder43sheet5C34B027B 1K
R409 alualuadder41adder43sheet5C34B00DA alualuadder41adder43sheet5C34B00DAorB 10K
R410 aluAdderB3in alualuadder41adder43sheet5C34B00DAorB 10K
Q169 alualuadder41adder43sheet5C34B027B alualuadder41adder43sheet5C34B00DAorB 0 NPN
R414 aluVcc alualuadder41adder43sheet5C34B047A 1K
R412 alualuadder41adder43sheet5C34B027A alualuadder41adder43sheet5C34B027AorB 10K
R413 alualuadder41adder43sheet5C34B027B alualuadder41adder43sheet5C34B027AorB 10K
Q170 alualuadder41adder43sheet5C34B047A alualuadder41adder43sheet5C34B027AorB 0 NPN
R417 aluVcc alualuadder41adder43sheet5C34B049A 1K
R415 alualuadder41adder43sheet5C34B047A alualuadder41adder43sheet5C34B047AorB 10K
R416 alualuadder41adder43Cin alualuadder41adder43sheet5C34B047AorB 10K
Q171 alualuadder41adder43sheet5C34B049A alualuadder41adder43sheet5C34B047AorB 0 NPN
R420 aluVcc alualuadder41adder43sheet5C34B04AA 1K
R418 alualuadder41adder43sheet5C34B047A alualuadder41adder43sheet5C34B048AorB 10K
R419 alualuadder41adder43sheet5C34B049A alualuadder41adder43sheet5C34B048AorB 10K
Q172 alualuadder41adder43sheet5C34B04AA alualuadder41adder43sheet5C34B048AorB 0 NPN
R423 aluVcc alualuadder41adder43sheet5C34B04AB 1K
R421 alualuadder41adder43sheet5C34B049A alualuadder41adder43sheet5C34B049AorB 10K
R422 alualuadder41adder43Cin alualuadder41adder43sheet5C34B049AorB 10K
Q173 alualuadder41adder43sheet5C34B04AB alualuadder41adder43sheet5C34B049AorB 0 NPN
R426 aluVcc aluAdderS3 1K
R424 alualuadder41adder43sheet5C34B04AA alualuadder41adder43sheet5C34B04AAorB 10K
R425 alualuadder41adder43sheet5C34B04AB alualuadder41adder43sheet5C34B04AAorB 10K
Q174 aluAdderS3 alualuadder41adder43sheet5C34B04AAorB 0 NPN
R429 aluVcc alualuadder41adder44Cin 1K
R427 alualuadder41adder43sheet5C34B049A alualuadder41adder43sheet5C34B0CDAorB 10K
R428 alualuadder41adder43sheet5C34B00DA alualuadder41adder43sheet5C34B0CDAorB 10K
Q175 alualuadder41adder44Cin alualuadder41adder43sheet5C34B0CDAorB 0 NPN
R432 aluVcc alualuadder41adder44sheet5C34B00DA 1K
R430 A4in alualuadder41adder44sheet5C34AF27AorB 10K
R431 aluAdderB4in alualuadder41adder44sheet5C34AF27AorB 10K
Q176 alualuadder41adder44sheet5C34B00DA alualuadder41adder44sheet5C34AF27AorB 0 NPN
R435 aluVcc alualuadder41adder44sheet5C34B027A 1K
R433 A4in alualuadder41adder44sheet5C34AFF9AorB 10K
R434 alualuadder41adder44sheet5C34B00DA alualuadder41adder44sheet5C34AFF9AorB 10K
Q177 alualuadder41adder44sheet5C34B027A alualuadder41adder44sheet5C34AFF9AorB 0 NPN
R438 aluVcc alualuadder41adder44sheet5C34B027B 1K
R436 alualuadder41adder44sheet5C34B00DA alualuadder41adder44sheet5C34B00DAorB 10K
R437 aluAdderB4in alualuadder41adder44sheet5C34B00DAorB 10K
Q178 alualuadder41adder44sheet5C34B027B alualuadder41adder44sheet5C34B00DAorB 0 NPN
R441 aluVcc alualuadder41adder44sheet5C34B047A 1K
R439 alualuadder41adder44sheet5C34B027A alualuadder41adder44sheet5C34B027AorB 10K
R440 alualuadder41adder44sheet5C34B027B alualuadder41adder44sheet5C34B027AorB 10K
Q179 alualuadder41adder44sheet5C34B047A alualuadder41adder44sheet5C34B027AorB 0 NPN
R444 aluVcc alualuadder41adder44sheet5C34B049A 1K
R442 alualuadder41adder44sheet5C34B047A alualuadder41adder44sheet5C34B047AorB 10K
R443 alualuadder41adder44Cin alualuadder41adder44sheet5C34B047AorB 10K
Q180 alualuadder41adder44sheet5C34B049A alualuadder41adder44sheet5C34B047AorB 0 NPN
R447 aluVcc alualuadder41adder44sheet5C34B04AA 1K
R445 alualuadder41adder44sheet5C34B047A alualuadder41adder44sheet5C34B048AorB 10K
R446 alualuadder41adder44sheet5C34B049A alualuadder41adder44sheet5C34B048AorB 10K
Q181 alualuadder41adder44sheet5C34B04AA alualuadder41adder44sheet5C34B048AorB 0 NPN
R450 aluVcc alualuadder41adder44sheet5C34B04AB 1K
R448 alualuadder41adder44sheet5C34B049A alualuadder41adder44sheet5C34B049AorB 10K
R449 alualuadder41adder44Cin alualuadder41adder44sheet5C34B049AorB 10K
Q182 alualuadder41adder44sheet5C34B04AB alualuadder41adder44sheet5C34B049AorB 0 NPN
R453 aluVcc aluAdderS4 1K
R451 alualuadder41adder44sheet5C34B04AA alualuadder41adder44sheet5C34B04AAorB 10K
R452 alualuadder41adder44sheet5C34B04AB alualuadder41adder44sheet5C34B04AAorB 10K
Q183 aluAdderS4 alualuadder41adder44sheet5C34B04AAorB 0 NPN
R456 aluVcc aluCout 1K
R454 alualuadder41adder44sheet5C34B049A alualuadder41adder44sheet5C34B0CDAorB 10K
R455 alualuadder41adder44sheet5C34B00DA alualuadder41adder44sheet5C34B0CDAorB 10K
Q184 aluCout alualuadder41adder44sheet5C34B0CDAorB 0 NPN
R459 aluVcc aluAdderB1in 1K
R457 alualuand41gateand42and1sheet5C364DB7A alualuand41gateand42and1sheet5C364DB7AorB 10K
R458 alualuand41gateand42and1sheet5C364DB7B alualuand41gateand42and1sheet5C364DB7AorB 10K
Q185 aluAdderB1in alualuand41gateand42and1sheet5C364DB7AorB 0 NPN
R461 aluVcc alualuand41gateand42and1sheet5C364DB7A 1K
R460 alualuand41A1 alualuand41gateand42and1Sheet5C3654CCQr 10K
Q186 alualuand41gateand42and1sheet5C364DB7A alualuand41gateand42and1Sheet5C3654CCQr 0 NPN
R463 aluVcc alualuand41gateand42and1sheet5C364DB7B 1K
R462 alualuand41B1 alualuand41gateand42and1sheet5C366192Qr 10K
Q187 alualuand41gateand42and1sheet5C364DB7B alualuand41gateand42and1sheet5C366192Qr 0 NPN
R466 aluVcc aluAdderB2in 1K
R464 alualuand41gateand42and2sheet5C364DB7A alualuand41gateand42and2sheet5C364DB7AorB 10K
R465 alualuand41gateand42and2sheet5C364DB7B alualuand41gateand42and2sheet5C364DB7AorB 10K
Q188 aluAdderB2in alualuand41gateand42and2sheet5C364DB7AorB 0 NPN
R468 aluVcc alualuand41gateand42and2sheet5C364DB7A 1K
R467 alualuand41A2 alualuand41gateand42and2Sheet5C3654CCQr 10K
Q189 alualuand41gateand42and2sheet5C364DB7A alualuand41gateand42and2Sheet5C3654CCQr 0 NPN
R470 aluVcc alualuand41gateand42and2sheet5C364DB7B 1K
R469 alualuand41B2 alualuand41gateand42and2sheet5C366192Qr 10K
Q190 alualuand41gateand42and2sheet5C364DB7B alualuand41gateand42and2sheet5C366192Qr 0 NPN
R473 aluVcc aluAdderB3in 1K
R471 alualuand41gateand42and3sheet5C364DB7A alualuand41gateand42and3sheet5C364DB7AorB 10K
R472 alualuand41gateand42and3sheet5C364DB7B alualuand41gateand42and3sheet5C364DB7AorB 10K
Q191 aluAdderB3in alualuand41gateand42and3sheet5C364DB7AorB 0 NPN
R475 aluVcc alualuand41gateand42and3sheet5C364DB7A 1K
R474 alualuand41A3 alualuand41gateand42and3Sheet5C3654CCQr 10K
Q192 alualuand41gateand42and3sheet5C364DB7A alualuand41gateand42and3Sheet5C3654CCQr 0 NPN
R477 aluVcc alualuand41gateand42and3sheet5C364DB7B 1K
R476 alualuand41B3 alualuand41gateand42and3sheet5C366192Qr 10K
Q193 alualuand41gateand42and3sheet5C364DB7B alualuand41gateand42and3sheet5C366192Qr 0 NPN
R480 aluVcc aluAdderB4in 1K
R478 alualuand41gateand42and4sheet5C364DB7A alualuand41gateand42and4sheet5C364DB7AorB 10K
R479 alualuand41gateand42and4sheet5C364DB7B alualuand41gateand42and4sheet5C364DB7AorB 10K
Q194 aluAdderB4in alualuand41gateand42and4sheet5C364DB7AorB 0 NPN
R482 aluVcc alualuand41gateand42and4sheet5C364DB7A 1K
R481 alualuand41A4 alualuand41gateand42and4Sheet5C3654CCQr 10K
Q195 alualuand41gateand42and4sheet5C364DB7A alualuand41gateand42and4Sheet5C3654CCQr 0 NPN
R484 aluVcc alualuand41gateand42and4sheet5C364DB7B 1K
R483 alualuand41B4 alualuand41gateand42and4sheet5C366192Qr 10K
Q196 alualuand41gateand42and4sheet5C364DB7B alualuand41gateand42and4sheet5C366192Qr 0 NPN
R486 aluVcc alualureplicate141A 1K
R485 S5 alualunot1Qr 10K
Q197 alualureplicate141A alualunot1Qr 0 NPN
.end
