.title KiCad schematic
V1 /nor-2/Vcc 0 dc 5
V2 /Ain 0 dc 5
V3 /Bin 0 dc 5
R3 /nor-2/Vcc /Q 1K
R1 /Ain /nor-2/AorB 10K
R2 /Bin /nor-2/AorB 10K
Q1 /Q /nor-2/AorB 0 NPN
.end
