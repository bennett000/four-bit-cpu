.title KiCad schematic
.op
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V1 multiplexer421Vcc 0 dc 5
V2 A1in 0 dc 5
V3 A2in 0 dc 0
V4 A3in 0 dc 5
V5 A4in 0 dc 0
V9 B4in 0 dc 0
V8 B3in 0 dc 5
V7 B2in 0 dc 5
V6 B1in 0 dc 0
V10 SelIn 0 dc 5
R2 multiplexer421Vcc multiplexer421Z1 1K
R1 multiplexer421multiplexer421mux1211mux21or1ornor1Q multiplexer421multiplexer421mux1211mux21or1ornot1Qr 10K
Q1 multiplexer421Z1 multiplexer421multiplexer421mux1211mux21or1ornot1Qr 0 NPN
R5 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21or1ornor1Q 1K
R3 multiplexer421multiplexer421mux1211mux21or1A multiplexer421multiplexer421mux1211mux21or1ornor1AorB 10K
R4 multiplexer421multiplexer421mux1211mux21or1B multiplexer421multiplexer421mux1211mux21or1ornor1AorB 10K
Q2 multiplexer421multiplexer421mux1211mux21or1ornor1Q multiplexer421multiplexer421mux1211mux21or1ornor1AorB 0 NPN
R8 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21or1A 1K
R6 multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
R7 multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7AorB 10K
Q3 multiplexer421multiplexer421mux1211mux21or1A multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7AorB 0 NPN
R10 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7A 1K
R9 A1in multiplexer421multiplexer421mux1211mux21and1Sheet5C3654CCQr 10K
Q4 multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1211mux21and1Sheet5C3654CCQr 0 NPN
R12 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7B 1K
R11 multiplexer421multiplexer421mux1211mux21and1B multiplexer421multiplexer421mux1211mux21and1sheet5C366192Qr 10K
Q5 multiplexer421multiplexer421mux1211mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1211mux21and1sheet5C366192Qr 0 NPN
R15 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21or1B 1K
R13 multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
R14 multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7AorB 10K
Q6 multiplexer421multiplexer421mux1211mux21or1B multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7AorB 0 NPN
R17 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7A 1K
R16 SelIn multiplexer421multiplexer421mux1211mux21and2Sheet5C3654CCQr 10K
Q7 multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1211mux21and2Sheet5C3654CCQr 0 NPN
R19 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7B 1K
R18 B1in multiplexer421multiplexer421mux1211mux21and2sheet5C366192Qr 10K
Q8 multiplexer421multiplexer421mux1211mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1211mux21and2sheet5C366192Qr 0 NPN
R21 multiplexer421Vcc multiplexer421multiplexer421mux1211mux21and1B 1K
R20 SelIn multiplexer421multiplexer421mux1211mux21not1Qr 10K
Q9 multiplexer421multiplexer421mux1211mux21and1B multiplexer421multiplexer421mux1211mux21not1Qr 0 NPN
R23 multiplexer421Vcc multiplexer421Z2 1K
R22 multiplexer421multiplexer421mux1212mux21or1ornor1Q multiplexer421multiplexer421mux1212mux21or1ornot1Qr 10K
Q10 multiplexer421Z2 multiplexer421multiplexer421mux1212mux21or1ornot1Qr 0 NPN
R26 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21or1ornor1Q 1K
R24 multiplexer421multiplexer421mux1212mux21or1A multiplexer421multiplexer421mux1212mux21or1ornor1AorB 10K
R25 multiplexer421multiplexer421mux1212mux21or1B multiplexer421multiplexer421mux1212mux21or1ornor1AorB 10K
Q11 multiplexer421multiplexer421mux1212mux21or1ornor1Q multiplexer421multiplexer421mux1212mux21or1ornor1AorB 0 NPN
R29 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21or1A 1K
R27 multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
R28 multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7AorB 10K
Q12 multiplexer421multiplexer421mux1212mux21or1A multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7AorB 0 NPN
R31 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7A 1K
R30 A2in multiplexer421multiplexer421mux1212mux21and1Sheet5C3654CCQr 10K
Q13 multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1212mux21and1Sheet5C3654CCQr 0 NPN
R33 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7B 1K
R32 multiplexer421multiplexer421mux1212mux21and1B multiplexer421multiplexer421mux1212mux21and1sheet5C366192Qr 10K
Q14 multiplexer421multiplexer421mux1212mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1212mux21and1sheet5C366192Qr 0 NPN
R36 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21or1B 1K
R34 multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
R35 multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7AorB 10K
Q15 multiplexer421multiplexer421mux1212mux21or1B multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7AorB 0 NPN
R38 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7A 1K
R37 SelIn multiplexer421multiplexer421mux1212mux21and2Sheet5C3654CCQr 10K
Q16 multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1212mux21and2Sheet5C3654CCQr 0 NPN
R40 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7B 1K
R39 B2in multiplexer421multiplexer421mux1212mux21and2sheet5C366192Qr 10K
Q17 multiplexer421multiplexer421mux1212mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1212mux21and2sheet5C366192Qr 0 NPN
R42 multiplexer421Vcc multiplexer421multiplexer421mux1212mux21and1B 1K
R41 SelIn multiplexer421multiplexer421mux1212mux21not1Qr 10K
Q18 multiplexer421multiplexer421mux1212mux21and1B multiplexer421multiplexer421mux1212mux21not1Qr 0 NPN
R44 multiplexer421Vcc multiplexer421Z3 1K
R43 multiplexer421multiplexer421mux1213mux21or1ornor1Q multiplexer421multiplexer421mux1213mux21or1ornot1Qr 10K
Q19 multiplexer421Z3 multiplexer421multiplexer421mux1213mux21or1ornot1Qr 0 NPN
R47 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21or1ornor1Q 1K
R45 multiplexer421multiplexer421mux1213mux21or1A multiplexer421multiplexer421mux1213mux21or1ornor1AorB 10K
R46 multiplexer421multiplexer421mux1213mux21or1B multiplexer421multiplexer421mux1213mux21or1ornor1AorB 10K
Q20 multiplexer421multiplexer421mux1213mux21or1ornor1Q multiplexer421multiplexer421mux1213mux21or1ornor1AorB 0 NPN
R50 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21or1A 1K
R48 multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
R49 multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7AorB 10K
Q21 multiplexer421multiplexer421mux1213mux21or1A multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7AorB 0 NPN
R52 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7A 1K
R51 A3in multiplexer421multiplexer421mux1213mux21and1Sheet5C3654CCQr 10K
Q22 multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1213mux21and1Sheet5C3654CCQr 0 NPN
R54 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7B 1K
R53 multiplexer421multiplexer421mux1213mux21and1B multiplexer421multiplexer421mux1213mux21and1sheet5C366192Qr 10K
Q23 multiplexer421multiplexer421mux1213mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1213mux21and1sheet5C366192Qr 0 NPN
R57 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21or1B 1K
R55 multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
R56 multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7AorB 10K
Q24 multiplexer421multiplexer421mux1213mux21or1B multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7AorB 0 NPN
R59 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7A 1K
R58 SelIn multiplexer421multiplexer421mux1213mux21and2Sheet5C3654CCQr 10K
Q25 multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1213mux21and2Sheet5C3654CCQr 0 NPN
R61 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7B 1K
R60 B3in multiplexer421multiplexer421mux1213mux21and2sheet5C366192Qr 10K
Q26 multiplexer421multiplexer421mux1213mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1213mux21and2sheet5C366192Qr 0 NPN
R63 multiplexer421Vcc multiplexer421multiplexer421mux1213mux21and1B 1K
R62 SelIn multiplexer421multiplexer421mux1213mux21not1Qr 10K
Q27 multiplexer421multiplexer421mux1213mux21and1B multiplexer421multiplexer421mux1213mux21not1Qr 0 NPN
R65 multiplexer421Vcc multiplexer421Z4 1K
R64 multiplexer421multiplexer421mux1214mux21or1ornor1Q multiplexer421multiplexer421mux1214mux21or1ornot1Qr 10K
Q28 multiplexer421Z4 multiplexer421multiplexer421mux1214mux21or1ornot1Qr 0 NPN
R68 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21or1ornor1Q 1K
R66 multiplexer421multiplexer421mux1214mux21or1A multiplexer421multiplexer421mux1214mux21or1ornor1AorB 10K
R67 multiplexer421multiplexer421mux1214mux21or1B multiplexer421multiplexer421mux1214mux21or1ornor1AorB 10K
Q29 multiplexer421multiplexer421mux1214mux21or1ornor1Q multiplexer421multiplexer421mux1214mux21or1ornor1AorB 0 NPN
R71 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21or1A 1K
R69 multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
R70 multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7AorB 10K
Q30 multiplexer421multiplexer421mux1214mux21or1A multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7AorB 0 NPN
R73 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7A 1K
R72 A4in multiplexer421multiplexer421mux1214mux21and1Sheet5C3654CCQr 10K
Q31 multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7A multiplexer421multiplexer421mux1214mux21and1Sheet5C3654CCQr 0 NPN
R75 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7B 1K
R74 multiplexer421multiplexer421mux1214mux21and1B multiplexer421multiplexer421mux1214mux21and1sheet5C366192Qr 10K
Q32 multiplexer421multiplexer421mux1214mux21and1sheet5C364DB7B multiplexer421multiplexer421mux1214mux21and1sheet5C366192Qr 0 NPN
R78 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21or1B 1K
R76 multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
R77 multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7AorB 10K
Q33 multiplexer421multiplexer421mux1214mux21or1B multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7AorB 0 NPN
R80 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7A 1K
R79 SelIn multiplexer421multiplexer421mux1214mux21and2Sheet5C3654CCQr 10K
Q34 multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7A multiplexer421multiplexer421mux1214mux21and2Sheet5C3654CCQr 0 NPN
R82 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7B 1K
R81 B4in multiplexer421multiplexer421mux1214mux21and2sheet5C366192Qr 10K
Q35 multiplexer421multiplexer421mux1214mux21and2sheet5C364DB7B multiplexer421multiplexer421mux1214mux21and2sheet5C366192Qr 0 NPN
R84 multiplexer421Vcc multiplexer421multiplexer421mux1214mux21and1B 1K
R83 SelIn multiplexer421multiplexer421mux1214mux21not1Qr 10K
Q36 multiplexer421multiplexer421mux1214mux21and1B multiplexer421multiplexer421mux1214mux21not1Qr 0 NPN
.end
