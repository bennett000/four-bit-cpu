.title KiCad schematic
.op
.model NPN npn (is=6.7e-15 bf=416.4 nf=1 vaf=74.03 ikf=0.06678 ise=6.7e-15 ne=1.259 br=0.7371 nr=1 rb=10 rc=1)
V1 /not/Q 0 dc 5
R2 /not/Q /not/NQ 1K
*R1 /not/Q /not/Qr 10K
Q1 /not/NQ /not/Qr 0 NPN
.end
