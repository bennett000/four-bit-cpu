.title KiCad schematic
V1 /nor-3/Vcc 0 dc 5
V2 /Ain 0 dc 5
V3 /Bin 0 dc 5
V4 /Cin 0 dc 5
R4 /nor-3/Vcc /nor-3/Q 1K
R1 /Ain /nor-3/AorBorC 10K
R2 /Bin /nor-3/AorBorC 10K
Q1 /nor-3/Q /nor-3/AorBorC 0 NPN
R3 /Cin /nor-3/AorBorC 10K
.end
